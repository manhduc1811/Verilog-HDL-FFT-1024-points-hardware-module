module ROM_256(
input clk,
input in_valid,
input rst_n,
output reg [23:0] w_r,
output reg [23:0] w_i,
output reg[1:0] state
);

reg valid;
reg [10:0] count,next_count;
reg [8:0] s_count,next_s_count;

always @(*) begin
    if(in_valid || valid)
    begin 
        next_count = count + 1;
        next_s_count = s_count;
    end
    else begin
        next_count = count;
        next_s_count = s_count;  
    end
    
    if (count<11'd256) 
        state = 2'd0;
    else if (count >= 11'd256 && s_count < 9'd256)begin
        state = 2'd1;
        next_s_count = s_count + 1;
    end
    else if (count >= 11'd256 && s_count >= 9'd256)begin
        state = 2'd2;
        next_s_count = s_count + 1;
    end

	case(s_count)
	9'd256: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 000000000000000000000000;
	 end
	9'd257: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111111101;
	 end
	9'd258: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111111010;
	 end
	9'd259: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110111;
	 end
	9'd260: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110011;
	 end
	9'd261: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110000;
	 end
	9'd262: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111101101;
	 end
	9'd263: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111101010;
	 end
	9'd264: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111100111;
	 end
	9'd265: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111100100;
	 end
	9'd266: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111100001;
	 end
	9'd267: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111011110;
	 end
	9'd268: begin 
	 w_r = 24'b 000000000000000011111101;
	 w_i = 24'b 111111111111111111011010;
	 end
	9'd269: begin 
	 w_r = 24'b 000000000000000011111101;
	 w_i = 24'b 111111111111111111010111;
	 end
	9'd270: begin 
	 w_r = 24'b 000000000000000011111100;
	 w_i = 24'b 111111111111111111010100;
	 end
	9'd271: begin 
	 w_r = 24'b 000000000000000011111100;
	 w_i = 24'b 111111111111111111010001;
	 end
	9'd272: begin 
	 w_r = 24'b 000000000000000011111011;
	 w_i = 24'b 111111111111111111001110;
	 end
	9'd273: begin 
	 w_r = 24'b 000000000000000011111010;
	 w_i = 24'b 111111111111111111001011;
	 end
	9'd274: begin 
	 w_r = 24'b 000000000000000011111010;
	 w_i = 24'b 111111111111111111001000;
	 end
	9'd275: begin 
	 w_r = 24'b 000000000000000011111001;
	 w_i = 24'b 111111111111111111000101;
	 end
	9'd276: begin 
	 w_r = 24'b 000000000000000011111000;
	 w_i = 24'b 111111111111111111000010;
	 end
	9'd277: begin 
	 w_r = 24'b 000000000000000011111000;
	 w_i = 24'b 111111111111111110111111;
	 end
	9'd278: begin 
	 w_r = 24'b 000000000000000011110111;
	 w_i = 24'b 111111111111111110111100;
	 end
	9'd279: begin 
	 w_r = 24'b 000000000000000011110110;
	 w_i = 24'b 111111111111111110111001;
	 end
	9'd280: begin 
	 w_r = 24'b 000000000000000011110101;
	 w_i = 24'b 111111111111111110110110;
	 end
	9'd281: begin 
	 w_r = 24'b 000000000000000011110100;
	 w_i = 24'b 111111111111111110110011;
	 end
	9'd282: begin 
	 w_r = 24'b 000000000000000011110011;
	 w_i = 24'b 111111111111111110110000;
	 end
	9'd283: begin 
	 w_r = 24'b 000000000000000011110010;
	 w_i = 24'b 111111111111111110101101;
	 end
	9'd284: begin 
	 w_r = 24'b 000000000000000011110001;
	 w_i = 24'b 111111111111111110101010;
	 end
	9'd285: begin 
	 w_r = 24'b 000000000000000011110000;
	 w_i = 24'b 111111111111111110100111;
	 end
	9'd286: begin 
	 w_r = 24'b 000000000000000011101111;
	 w_i = 24'b 111111111111111110100100;
	 end
	9'd287: begin 
	 w_r = 24'b 000000000000000011101110;
	 w_i = 24'b 111111111111111110100001;
	 end
	9'd288: begin 
	 w_r = 24'b 000000000000000011101101;
	 w_i = 24'b 111111111111111110011110;
	 end
	9'd289: begin 
	 w_r = 24'b 000000000000000011101011;
	 w_i = 24'b 111111111111111110011011;
	 end
	9'd290: begin 
	 w_r = 24'b 000000000000000011101010;
	 w_i = 24'b 111111111111111110011000;
	 end
	9'd291: begin 
	 w_r = 24'b 000000000000000011101001;
	 w_i = 24'b 111111111111111110010101;
	 end
	9'd292: begin 
	 w_r = 24'b 000000000000000011100111;
	 w_i = 24'b 111111111111111110010011;
	 end
	9'd293: begin 
	 w_r = 24'b 000000000000000011100110;
	 w_i = 24'b 111111111111111110010000;
	 end
	9'd294: begin 
	 w_r = 24'b 000000000000000011100101;
	 w_i = 24'b 111111111111111110001101;
	 end
	9'd295: begin 
	 w_r = 24'b 000000000000000011100011;
	 w_i = 24'b 111111111111111110001010;
	 end
	9'd296: begin 
	 w_r = 24'b 000000000000000011100010;
	 w_i = 24'b 111111111111111110000111;
	 end
	9'd297: begin 
	 w_r = 24'b 000000000000000011100000;
	 w_i = 24'b 111111111111111110000101;
	 end
	9'd298: begin 
	 w_r = 24'b 000000000000000011011111;
	 w_i = 24'b 111111111111111110000010;
	 end
	9'd299: begin 
	 w_r = 24'b 000000000000000011011101;
	 w_i = 24'b 111111111111111101111111;
	 end
	9'd300: begin 
	 w_r = 24'b 000000000000000011011100;
	 w_i = 24'b 111111111111111101111100;
	 end
	9'd301: begin 
	 w_r = 24'b 000000000000000011011010;
	 w_i = 24'b 111111111111111101111010;
	 end
	9'd302: begin 
	 w_r = 24'b 000000000000000011011000;
	 w_i = 24'b 111111111111111101110111;
	 end
	9'd303: begin 
	 w_r = 24'b 000000000000000011010111;
	 w_i = 24'b 111111111111111101110100;
	 end
	9'd304: begin 
	 w_r = 24'b 000000000000000011010101;
	 w_i = 24'b 111111111111111101110010;
	 end
	9'd305: begin 
	 w_r = 24'b 000000000000000011010011;
	 w_i = 24'b 111111111111111101101111;
	 end
	9'd306: begin 
	 w_r = 24'b 000000000000000011010001;
	 w_i = 24'b 111111111111111101101101;
	 end
	9'd307: begin 
	 w_r = 24'b 000000000000000011001111;
	 w_i = 24'b 111111111111111101101010;
	 end
	9'd308: begin 
	 w_r = 24'b 000000000000000011001110;
	 w_i = 24'b 111111111111111101101000;
	 end
	9'd309: begin 
	 w_r = 24'b 000000000000000011001100;
	 w_i = 24'b 111111111111111101100101;
	 end
	9'd310: begin 
	 w_r = 24'b 000000000000000011001010;
	 w_i = 24'b 111111111111111101100011;
	 end
	9'd311: begin 
	 w_r = 24'b 000000000000000011001000;
	 w_i = 24'b 111111111111111101100000;
	 end
	9'd312: begin 
	 w_r = 24'b 000000000000000011000110;
	 w_i = 24'b 111111111111111101011110;
	 end
	9'd313: begin 
	 w_r = 24'b 000000000000000011000100;
	 w_i = 24'b 111111111111111101011011;
	 end
	9'd314: begin 
	 w_r = 24'b 000000000000000011000010;
	 w_i = 24'b 111111111111111101011001;
	 end
	9'd315: begin 
	 w_r = 24'b 000000000000000011000000;
	 w_i = 24'b 111111111111111101010110;
	 end
	9'd316: begin 
	 w_r = 24'b 000000000000000010111110;
	 w_i = 24'b 111111111111111101010100;
	 end
	9'd317: begin 
	 w_r = 24'b 000000000000000010111100;
	 w_i = 24'b 111111111111111101010010;
	 end
	9'd318: begin 
	 w_r = 24'b 000000000000000010111001;
	 w_i = 24'b 111111111111111101001111;
	 end
	9'd319: begin 
	 w_r = 24'b 000000000000000010110111;
	 w_i = 24'b 111111111111111101001101;
	 end
	9'd320: begin 
	 w_r = 24'b 000000000000000010110101;
	 w_i = 24'b 111111111111111101001011;
	 end
	9'd321: begin 
	 w_r = 24'b 000000000000000010110011;
	 w_i = 24'b 111111111111111101001001;
	 end
	9'd322: begin 
	 w_r = 24'b 000000000000000010110001;
	 w_i = 24'b 111111111111111101000111;
	 end
	9'd323: begin 
	 w_r = 24'b 000000000000000010101110;
	 w_i = 24'b 111111111111111101000100;
	 end
	9'd324: begin 
	 w_r = 24'b 000000000000000010101100;
	 w_i = 24'b 111111111111111101000010;
	 end
	9'd325: begin 
	 w_r = 24'b 000000000000000010101010;
	 w_i = 24'b 111111111111111101000000;
	 end
	9'd326: begin 
	 w_r = 24'b 000000000000000010100111;
	 w_i = 24'b 111111111111111100111110;
	 end
	9'd327: begin 
	 w_r = 24'b 000000000000000010100101;
	 w_i = 24'b 111111111111111100111100;
	 end
	9'd328: begin 
	 w_r = 24'b 000000000000000010100010;
	 w_i = 24'b 111111111111111100111010;
	 end
	9'd329: begin 
	 w_r = 24'b 000000000000000010100000;
	 w_i = 24'b 111111111111111100111000;
	 end
	9'd330: begin 
	 w_r = 24'b 000000000000000010011101;
	 w_i = 24'b 111111111111111100110110;
	 end
	9'd331: begin 
	 w_r = 24'b 000000000000000010011011;
	 w_i = 24'b 111111111111111100110100;
	 end
	9'd332: begin 
	 w_r = 24'b 000000000000000010011000;
	 w_i = 24'b 111111111111111100110010;
	 end
	9'd333: begin 
	 w_r = 24'b 000000000000000010010110;
	 w_i = 24'b 111111111111111100110001;
	 end
	9'd334: begin 
	 w_r = 24'b 000000000000000010010011;
	 w_i = 24'b 111111111111111100101111;
	 end
	9'd335: begin 
	 w_r = 24'b 000000000000000010010001;
	 w_i = 24'b 111111111111111100101101;
	 end
	9'd336: begin 
	 w_r = 24'b 000000000000000010001110;
	 w_i = 24'b 111111111111111100101011;
	 end
	9'd337: begin 
	 w_r = 24'b 000000000000000010001100;
	 w_i = 24'b 111111111111111100101001;
	 end
	9'd338: begin 
	 w_r = 24'b 000000000000000010001001;
	 w_i = 24'b 111111111111111100101000;
	 end
	9'd339: begin 
	 w_r = 24'b 000000000000000010000110;
	 w_i = 24'b 111111111111111100100110;
	 end
	9'd340: begin 
	 w_r = 24'b 000000000000000010000100;
	 w_i = 24'b 111111111111111100100100;
	 end
	9'd341: begin 
	 w_r = 24'b 000000000000000010000001;
	 w_i = 24'b 111111111111111100100011;
	 end
	9'd342: begin 
	 w_r = 24'b 000000000000000001111110;
	 w_i = 24'b 111111111111111100100001;
	 end
	9'd343: begin 
	 w_r = 24'b 000000000000000001111011;
	 w_i = 24'b 111111111111111100100000;
	 end
	9'd344: begin 
	 w_r = 24'b 000000000000000001111001;
	 w_i = 24'b 111111111111111100011110;
	 end
	9'd345: begin 
	 w_r = 24'b 000000000000000001110110;
	 w_i = 24'b 111111111111111100011101;
	 end
	9'd346: begin 
	 w_r = 24'b 000000000000000001110011;
	 w_i = 24'b 111111111111111100011011;
	 end
	9'd347: begin 
	 w_r = 24'b 000000000000000001110000;
	 w_i = 24'b 111111111111111100011010;
	 end
	9'd348: begin 
	 w_r = 24'b 000000000000000001101101;
	 w_i = 24'b 111111111111111100011001;
	 end
	9'd349: begin 
	 w_r = 24'b 000000000000000001101011;
	 w_i = 24'b 111111111111111100010111;
	 end
	9'd350: begin 
	 w_r = 24'b 000000000000000001101000;
	 w_i = 24'b 111111111111111100010110;
	 end
	9'd351: begin 
	 w_r = 24'b 000000000000000001100101;
	 w_i = 24'b 111111111111111100010101;
	 end
	9'd352: begin 
	 w_r = 24'b 000000000000000001100010;
	 w_i = 24'b 111111111111111100010011;
	 end
	9'd353: begin 
	 w_r = 24'b 000000000000000001011111;
	 w_i = 24'b 111111111111111100010010;
	 end
	9'd354: begin 
	 w_r = 24'b 000000000000000001011100;
	 w_i = 24'b 111111111111111100010001;
	 end
	9'd355: begin 
	 w_r = 24'b 000000000000000001011001;
	 w_i = 24'b 111111111111111100010000;
	 end
	9'd356: begin 
	 w_r = 24'b 000000000000000001010110;
	 w_i = 24'b 111111111111111100001111;
	 end
	9'd357: begin 
	 w_r = 24'b 000000000000000001010011;
	 w_i = 24'b 111111111111111100001110;
	 end
	9'd358: begin 
	 w_r = 24'b 000000000000000001010000;
	 w_i = 24'b 111111111111111100001101;
	 end
	9'd359: begin 
	 w_r = 24'b 000000000000000001001101;
	 w_i = 24'b 111111111111111100001100;
	 end
	9'd360: begin 
	 w_r = 24'b 000000000000000001001010;
	 w_i = 24'b 111111111111111100001011;
	 end
	9'd361: begin 
	 w_r = 24'b 000000000000000001000111;
	 w_i = 24'b 111111111111111100001010;
	 end
	9'd362: begin 
	 w_r = 24'b 000000000000000001000100;
	 w_i = 24'b 111111111111111100001001;
	 end
	9'd363: begin 
	 w_r = 24'b 000000000000000001000001;
	 w_i = 24'b 111111111111111100001000;
	 end
	9'd364: begin 
	 w_r = 24'b 000000000000000000111110;
	 w_i = 24'b 111111111111111100001000;
	 end
	9'd365: begin 
	 w_r = 24'b 000000000000000000111011;
	 w_i = 24'b 111111111111111100000111;
	 end
	9'd366: begin 
	 w_r = 24'b 000000000000000000111000;
	 w_i = 24'b 111111111111111100000110;
	 end
	9'd367: begin 
	 w_r = 24'b 000000000000000000110101;
	 w_i = 24'b 111111111111111100000110;
	 end
	9'd368: begin 
	 w_r = 24'b 000000000000000000110010;
	 w_i = 24'b 111111111111111100000101;
	 end
	9'd369: begin 
	 w_r = 24'b 000000000000000000101111;
	 w_i = 24'b 111111111111111100000100;
	 end
	9'd370: begin 
	 w_r = 24'b 000000000000000000101100;
	 w_i = 24'b 111111111111111100000100;
	 end
	9'd371: begin 
	 w_r = 24'b 000000000000000000101001;
	 w_i = 24'b 111111111111111100000011;
	 end
	9'd372: begin 
	 w_r = 24'b 000000000000000000100110;
	 w_i = 24'b 111111111111111100000011;
	 end
	9'd373: begin 
	 w_r = 24'b 000000000000000000100010;
	 w_i = 24'b 111111111111111100000010;
	 end
	9'd374: begin 
	 w_r = 24'b 000000000000000000011111;
	 w_i = 24'b 111111111111111100000010;
	 end
	9'd375: begin 
	 w_r = 24'b 000000000000000000011100;
	 w_i = 24'b 111111111111111100000010;
	 end
	9'd376: begin 
	 w_r = 24'b 000000000000000000011001;
	 w_i = 24'b 111111111111111100000001;
	 end
	9'd377: begin 
	 w_r = 24'b 000000000000000000010110;
	 w_i = 24'b 111111111111111100000001;
	 end
	9'd378: begin 
	 w_r = 24'b 000000000000000000010011;
	 w_i = 24'b 111111111111111100000001;
	 end
	9'd379: begin 
	 w_r = 24'b 000000000000000000010000;
	 w_i = 24'b 111111111111111100000000;
	 end
	9'd380: begin 
	 w_r = 24'b 000000000000000000001101;
	 w_i = 24'b 111111111111111100000000;
	 end
	9'd381: begin 
	 w_r = 24'b 000000000000000000001001;
	 w_i = 24'b 111111111111111100000000;
	 end
	9'd382: begin 
	 w_r = 24'b 000000000000000000000110;
	 w_i = 24'b 111111111111111100000000;
	 end
	9'd383: begin 
	 w_r = 24'b 000000000000000000000011;
	 w_i = 24'b 111111111111111100000000;
	 end
	9'd384: begin 
	 w_r = 24'b 000000000000000000000000;
	 w_i = 24'b 111111111111111100000000;
	 end
	9'd385: begin 
	 w_r = 24'b 111111111111111111111101;
	 w_i = 24'b 111111111111111100000000;
	 end
	9'd386: begin 
	 w_r = 24'b 111111111111111111111010;
	 w_i = 24'b 111111111111111100000000;
	 end
	9'd387: begin 
	 w_r = 24'b 111111111111111111110111;
	 w_i = 24'b 111111111111111100000000;
	 end
	9'd388: begin 
	 w_r = 24'b 111111111111111111110011;
	 w_i = 24'b 111111111111111100000000;
	 end
	9'd389: begin 
	 w_r = 24'b 111111111111111111110000;
	 w_i = 24'b 111111111111111100000000;
	 end
	9'd390: begin 
	 w_r = 24'b 111111111111111111101101;
	 w_i = 24'b 111111111111111100000001;
	 end
	9'd391: begin 
	 w_r = 24'b 111111111111111111101010;
	 w_i = 24'b 111111111111111100000001;
	 end
	9'd392: begin 
	 w_r = 24'b 111111111111111111100111;
	 w_i = 24'b 111111111111111100000001;
	 end
	9'd393: begin 
	 w_r = 24'b 111111111111111111100100;
	 w_i = 24'b 111111111111111100000010;
	 end
	9'd394: begin 
	 w_r = 24'b 111111111111111111100001;
	 w_i = 24'b 111111111111111100000010;
	 end
	9'd395: begin 
	 w_r = 24'b 111111111111111111011110;
	 w_i = 24'b 111111111111111100000010;
	 end
	9'd396: begin 
	 w_r = 24'b 111111111111111111011010;
	 w_i = 24'b 111111111111111100000011;
	 end
	9'd397: begin 
	 w_r = 24'b 111111111111111111010111;
	 w_i = 24'b 111111111111111100000011;
	 end
	9'd398: begin 
	 w_r = 24'b 111111111111111111010100;
	 w_i = 24'b 111111111111111100000100;
	 end
	9'd399: begin 
	 w_r = 24'b 111111111111111111010001;
	 w_i = 24'b 111111111111111100000100;
	 end
	9'd400: begin 
	 w_r = 24'b 111111111111111111001110;
	 w_i = 24'b 111111111111111100000101;
	 end
	9'd401: begin 
	 w_r = 24'b 111111111111111111001011;
	 w_i = 24'b 111111111111111100000110;
	 end
	9'd402: begin 
	 w_r = 24'b 111111111111111111001000;
	 w_i = 24'b 111111111111111100000110;
	 end
	9'd403: begin 
	 w_r = 24'b 111111111111111111000101;
	 w_i = 24'b 111111111111111100000111;
	 end
	9'd404: begin 
	 w_r = 24'b 111111111111111111000010;
	 w_i = 24'b 111111111111111100001000;
	 end
	9'd405: begin 
	 w_r = 24'b 111111111111111110111111;
	 w_i = 24'b 111111111111111100001000;
	 end
	9'd406: begin 
	 w_r = 24'b 111111111111111110111100;
	 w_i = 24'b 111111111111111100001001;
	 end
	9'd407: begin 
	 w_r = 24'b 111111111111111110111001;
	 w_i = 24'b 111111111111111100001010;
	 end
	9'd408: begin 
	 w_r = 24'b 111111111111111110110110;
	 w_i = 24'b 111111111111111100001011;
	 end
	9'd409: begin 
	 w_r = 24'b 111111111111111110110011;
	 w_i = 24'b 111111111111111100001100;
	 end
	9'd410: begin 
	 w_r = 24'b 111111111111111110110000;
	 w_i = 24'b 111111111111111100001101;
	 end
	9'd411: begin 
	 w_r = 24'b 111111111111111110101101;
	 w_i = 24'b 111111111111111100001110;
	 end
	9'd412: begin 
	 w_r = 24'b 111111111111111110101010;
	 w_i = 24'b 111111111111111100001111;
	 end
	9'd413: begin 
	 w_r = 24'b 111111111111111110100111;
	 w_i = 24'b 111111111111111100010000;
	 end
	9'd414: begin 
	 w_r = 24'b 111111111111111110100100;
	 w_i = 24'b 111111111111111100010001;
	 end
	9'd415: begin 
	 w_r = 24'b 111111111111111110100001;
	 w_i = 24'b 111111111111111100010010;
	 end
	9'd416: begin 
	 w_r = 24'b 111111111111111110011110;
	 w_i = 24'b 111111111111111100010011;
	 end
	9'd417: begin 
	 w_r = 24'b 111111111111111110011011;
	 w_i = 24'b 111111111111111100010101;
	 end
	9'd418: begin 
	 w_r = 24'b 111111111111111110011000;
	 w_i = 24'b 111111111111111100010110;
	 end
	9'd419: begin 
	 w_r = 24'b 111111111111111110010101;
	 w_i = 24'b 111111111111111100010111;
	 end
	9'd420: begin 
	 w_r = 24'b 111111111111111110010011;
	 w_i = 24'b 111111111111111100011001;
	 end
	9'd421: begin 
	 w_r = 24'b 111111111111111110010000;
	 w_i = 24'b 111111111111111100011010;
	 end
	9'd422: begin 
	 w_r = 24'b 111111111111111110001101;
	 w_i = 24'b 111111111111111100011011;
	 end
	9'd423: begin 
	 w_r = 24'b 111111111111111110001010;
	 w_i = 24'b 111111111111111100011101;
	 end
	9'd424: begin 
	 w_r = 24'b 111111111111111110000111;
	 w_i = 24'b 111111111111111100011110;
	 end
	9'd425: begin 
	 w_r = 24'b 111111111111111110000101;
	 w_i = 24'b 111111111111111100100000;
	 end
	9'd426: begin 
	 w_r = 24'b 111111111111111110000010;
	 w_i = 24'b 111111111111111100100001;
	 end
	9'd427: begin 
	 w_r = 24'b 111111111111111101111111;
	 w_i = 24'b 111111111111111100100011;
	 end
	9'd428: begin 
	 w_r = 24'b 111111111111111101111100;
	 w_i = 24'b 111111111111111100100100;
	 end
	9'd429: begin 
	 w_r = 24'b 111111111111111101111010;
	 w_i = 24'b 111111111111111100100110;
	 end
	9'd430: begin 
	 w_r = 24'b 111111111111111101110111;
	 w_i = 24'b 111111111111111100101000;
	 end
	9'd431: begin 
	 w_r = 24'b 111111111111111101110100;
	 w_i = 24'b 111111111111111100101001;
	 end
	9'd432: begin 
	 w_r = 24'b 111111111111111101110010;
	 w_i = 24'b 111111111111111100101011;
	 end
	9'd433: begin 
	 w_r = 24'b 111111111111111101101111;
	 w_i = 24'b 111111111111111100101101;
	 end
	9'd434: begin 
	 w_r = 24'b 111111111111111101101101;
	 w_i = 24'b 111111111111111100101111;
	 end
	9'd435: begin 
	 w_r = 24'b 111111111111111101101010;
	 w_i = 24'b 111111111111111100110001;
	 end
	9'd436: begin 
	 w_r = 24'b 111111111111111101101000;
	 w_i = 24'b 111111111111111100110010;
	 end
	9'd437: begin 
	 w_r = 24'b 111111111111111101100101;
	 w_i = 24'b 111111111111111100110100;
	 end
	9'd438: begin 
	 w_r = 24'b 111111111111111101100011;
	 w_i = 24'b 111111111111111100110110;
	 end
	9'd439: begin 
	 w_r = 24'b 111111111111111101100000;
	 w_i = 24'b 111111111111111100111000;
	 end
	9'd440: begin 
	 w_r = 24'b 111111111111111101011110;
	 w_i = 24'b 111111111111111100111010;
	 end
	9'd441: begin 
	 w_r = 24'b 111111111111111101011011;
	 w_i = 24'b 111111111111111100111100;
	 end
	9'd442: begin 
	 w_r = 24'b 111111111111111101011001;
	 w_i = 24'b 111111111111111100111110;
	 end
	9'd443: begin 
	 w_r = 24'b 111111111111111101010110;
	 w_i = 24'b 111111111111111101000000;
	 end
	9'd444: begin 
	 w_r = 24'b 111111111111111101010100;
	 w_i = 24'b 111111111111111101000010;
	 end
	9'd445: begin 
	 w_r = 24'b 111111111111111101010010;
	 w_i = 24'b 111111111111111101000100;
	 end
	9'd446: begin 
	 w_r = 24'b 111111111111111101001111;
	 w_i = 24'b 111111111111111101000111;
	 end
	9'd447: begin 
	 w_r = 24'b 111111111111111101001101;
	 w_i = 24'b 111111111111111101001001;
	 end
	9'd448: begin 
	 w_r = 24'b 111111111111111101001011;
	 w_i = 24'b 111111111111111101001011;
	 end
	9'd449: begin 
	 w_r = 24'b 111111111111111101001001;
	 w_i = 24'b 111111111111111101001101;
	 end
	9'd450: begin 
	 w_r = 24'b 111111111111111101000111;
	 w_i = 24'b 111111111111111101001111;
	 end
	9'd451: begin 
	 w_r = 24'b 111111111111111101000100;
	 w_i = 24'b 111111111111111101010010;
	 end
	9'd452: begin 
	 w_r = 24'b 111111111111111101000010;
	 w_i = 24'b 111111111111111101010100;
	 end
	9'd453: begin 
	 w_r = 24'b 111111111111111101000000;
	 w_i = 24'b 111111111111111101010110;
	 end
	9'd454: begin 
	 w_r = 24'b 111111111111111100111110;
	 w_i = 24'b 111111111111111101011001;
	 end
	9'd455: begin 
	 w_r = 24'b 111111111111111100111100;
	 w_i = 24'b 111111111111111101011011;
	 end
	9'd456: begin 
	 w_r = 24'b 111111111111111100111010;
	 w_i = 24'b 111111111111111101011110;
	 end
	9'd457: begin 
	 w_r = 24'b 111111111111111100111000;
	 w_i = 24'b 111111111111111101100000;
	 end
	9'd458: begin 
	 w_r = 24'b 111111111111111100110110;
	 w_i = 24'b 111111111111111101100011;
	 end
	9'd459: begin 
	 w_r = 24'b 111111111111111100110100;
	 w_i = 24'b 111111111111111101100101;
	 end
	9'd460: begin 
	 w_r = 24'b 111111111111111100110010;
	 w_i = 24'b 111111111111111101101000;
	 end
	9'd461: begin 
	 w_r = 24'b 111111111111111100110001;
	 w_i = 24'b 111111111111111101101010;
	 end
	9'd462: begin 
	 w_r = 24'b 111111111111111100101111;
	 w_i = 24'b 111111111111111101101101;
	 end
	9'd463: begin 
	 w_r = 24'b 111111111111111100101101;
	 w_i = 24'b 111111111111111101101111;
	 end
	9'd464: begin 
	 w_r = 24'b 111111111111111100101011;
	 w_i = 24'b 111111111111111101110010;
	 end
	9'd465: begin 
	 w_r = 24'b 111111111111111100101001;
	 w_i = 24'b 111111111111111101110100;
	 end
	9'd466: begin 
	 w_r = 24'b 111111111111111100101000;
	 w_i = 24'b 111111111111111101110111;
	 end
	9'd467: begin 
	 w_r = 24'b 111111111111111100100110;
	 w_i = 24'b 111111111111111101111010;
	 end
	9'd468: begin 
	 w_r = 24'b 111111111111111100100100;
	 w_i = 24'b 111111111111111101111100;
	 end
	9'd469: begin 
	 w_r = 24'b 111111111111111100100011;
	 w_i = 24'b 111111111111111101111111;
	 end
	9'd470: begin 
	 w_r = 24'b 111111111111111100100001;
	 w_i = 24'b 111111111111111110000010;
	 end
	9'd471: begin 
	 w_r = 24'b 111111111111111100100000;
	 w_i = 24'b 111111111111111110000101;
	 end
	9'd472: begin 
	 w_r = 24'b 111111111111111100011110;
	 w_i = 24'b 111111111111111110000111;
	 end
	9'd473: begin 
	 w_r = 24'b 111111111111111100011101;
	 w_i = 24'b 111111111111111110001010;
	 end
	9'd474: begin 
	 w_r = 24'b 111111111111111100011011;
	 w_i = 24'b 111111111111111110001101;
	 end
	9'd475: begin 
	 w_r = 24'b 111111111111111100011010;
	 w_i = 24'b 111111111111111110010000;
	 end
	9'd476: begin 
	 w_r = 24'b 111111111111111100011001;
	 w_i = 24'b 111111111111111110010011;
	 end
	9'd477: begin 
	 w_r = 24'b 111111111111111100010111;
	 w_i = 24'b 111111111111111110010101;
	 end
	9'd478: begin 
	 w_r = 24'b 111111111111111100010110;
	 w_i = 24'b 111111111111111110011000;
	 end
	9'd479: begin 
	 w_r = 24'b 111111111111111100010101;
	 w_i = 24'b 111111111111111110011011;
	 end
	9'd480: begin 
	 w_r = 24'b 111111111111111100010011;
	 w_i = 24'b 111111111111111110011110;
	 end
	9'd481: begin 
	 w_r = 24'b 111111111111111100010010;
	 w_i = 24'b 111111111111111110100001;
	 end
	9'd482: begin 
	 w_r = 24'b 111111111111111100010001;
	 w_i = 24'b 111111111111111110100100;
	 end
	9'd483: begin 
	 w_r = 24'b 111111111111111100010000;
	 w_i = 24'b 111111111111111110100111;
	 end
	9'd484: begin 
	 w_r = 24'b 111111111111111100001111;
	 w_i = 24'b 111111111111111110101010;
	 end
	9'd485: begin 
	 w_r = 24'b 111111111111111100001110;
	 w_i = 24'b 111111111111111110101101;
	 end
	9'd486: begin 
	 w_r = 24'b 111111111111111100001101;
	 w_i = 24'b 111111111111111110110000;
	 end
	9'd487: begin 
	 w_r = 24'b 111111111111111100001100;
	 w_i = 24'b 111111111111111110110011;
	 end
	9'd488: begin 
	 w_r = 24'b 111111111111111100001011;
	 w_i = 24'b 111111111111111110110110;
	 end
	9'd489: begin 
	 w_r = 24'b 111111111111111100001010;
	 w_i = 24'b 111111111111111110111001;
	 end
	9'd490: begin 
	 w_r = 24'b 111111111111111100001001;
	 w_i = 24'b 111111111111111110111100;
	 end
	9'd491: begin 
	 w_r = 24'b 111111111111111100001000;
	 w_i = 24'b 111111111111111110111111;
	 end
	9'd492: begin 
	 w_r = 24'b 111111111111111100001000;
	 w_i = 24'b 111111111111111111000010;
	 end
	9'd493: begin 
	 w_r = 24'b 111111111111111100000111;
	 w_i = 24'b 111111111111111111000101;
	 end
	9'd494: begin 
	 w_r = 24'b 111111111111111100000110;
	 w_i = 24'b 111111111111111111001000;
	 end
	9'd495: begin 
	 w_r = 24'b 111111111111111100000110;
	 w_i = 24'b 111111111111111111001011;
	 end
	9'd496: begin 
	 w_r = 24'b 111111111111111100000101;
	 w_i = 24'b 111111111111111111001110;
	 end
	9'd497: begin 
	 w_r = 24'b 111111111111111100000100;
	 w_i = 24'b 111111111111111111010001;
	 end
	9'd498: begin 
	 w_r = 24'b 111111111111111100000100;
	 w_i = 24'b 111111111111111111010100;
	 end
	9'd499: begin 
	 w_r = 24'b 111111111111111100000011;
	 w_i = 24'b 111111111111111111010111;
	 end
	9'd500: begin 
	 w_r = 24'b 111111111111111100000011;
	 w_i = 24'b 111111111111111111011010;
	 end
	9'd501: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111011110;
	 end
	9'd502: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111100001;
	 end
	9'd503: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111100100;
	 end
	9'd504: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111100111;
	 end
	9'd505: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111101010;
	 end
	9'd506: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111101101;
	 end
	9'd507: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110000;
	 end
	9'd508: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110011;
	 end
	9'd509: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110111;
	 end
	9'd510: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111111010;
	 end
	9'd511: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111111101;
	 end
	default: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 000000000000000000000000;
	 end
	endcase
end

always@(posedge clk or negedge rst_n)begin
    if(~rst_n)begin
        count <= 0;
        s_count <= 0;
    end
    else begin
        count <= next_count;
        s_count <= next_s_count;
    end
end
endmodule