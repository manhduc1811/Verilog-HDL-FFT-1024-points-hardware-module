module ROM_512(
input clk,
input in_valid,
input rst_n,
output reg [23:0] w_r,
output reg [23:0] w_i,
output reg[1:0] state
);

reg valid,next_valid;
reg [10:0] count,next_count;
always @(*) begin
    if(in_valid || valid)next_count = count + 1;
    else next_count = count;
    
    if (count<11'd512) 
        state = 2'd0;
    else if (count >= 11'd512 && count < 11'd1024)
        state = 2'd1;
    else if (count >= 11'd1024 && count < 11'd1536)
        state = 2'd2;
    else state = 2'd3;

	case(count)
	11'd1024: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 000000000000000000000000;
	 next_valid = 1'b1;
	 end
	11'd1025: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111111110;
	 next_valid = 1'b1;
	 end
	11'd1026: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111111101;
	 next_valid = 1'b1;
	 end
	11'd1027: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111111011;
	 next_valid = 1'b1;
	 end
	11'd1028: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111111010;
	 next_valid = 1'b1;
	 end
	11'd1029: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111111000;
	 next_valid = 1'b1;
	 end
	11'd1030: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110111;
	 next_valid = 1'b1;
	 end
	11'd1031: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110101;
	 next_valid = 1'b1;
	 end
	11'd1032: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110011;
	 next_valid = 1'b1;
	 end
	11'd1033: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110010;
	 next_valid = 1'b1;
	 end
	11'd1034: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110000;
	 next_valid = 1'b1;
	 end
	11'd1035: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111101111;
	 next_valid = 1'b1;
	 end
	11'd1036: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111101101;
	 next_valid = 1'b1;
	 end
	11'd1037: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111101100;
	 next_valid = 1'b1;
	 end
	11'd1038: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111101010;
	 next_valid = 1'b1;
	 end
	11'd1039: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111101000;
	 next_valid = 1'b1;
	 end
	11'd1040: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111100111;
	 next_valid = 1'b1;
	 end
	11'd1041: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111100101;
	 next_valid = 1'b1;
	 end
	11'd1042: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111100100;
	 next_valid = 1'b1;
	 end
	11'd1043: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111100010;
	 next_valid = 1'b1;
	 end
	11'd1044: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111100001;
	 next_valid = 1'b1;
	 end
	11'd1045: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111011111;
	 next_valid = 1'b1;
	 end
	11'd1046: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111011110;
	 next_valid = 1'b1;
	 end
	11'd1047: begin 
	 w_r = 24'b 000000000000000011111101;
	 w_i = 24'b 111111111111111111011100;
	 next_valid = 1'b1;
	 end
	11'd1048: begin 
	 w_r = 24'b 000000000000000011111101;
	 w_i = 24'b 111111111111111111011010;
	 next_valid = 1'b1;
	 end
	11'd1049: begin 
	 w_r = 24'b 000000000000000011111101;
	 w_i = 24'b 111111111111111111011001;
	 next_valid = 1'b1;
	 end
	11'd1050: begin 
	 w_r = 24'b 000000000000000011111101;
	 w_i = 24'b 111111111111111111010111;
	 next_valid = 1'b1;
	 end
	11'd1051: begin 
	 w_r = 24'b 000000000000000011111100;
	 w_i = 24'b 111111111111111111010110;
	 next_valid = 1'b1;
	 end
	11'd1052: begin 
	 w_r = 24'b 000000000000000011111100;
	 w_i = 24'b 111111111111111111010100;
	 next_valid = 1'b1;
	 end
	11'd1053: begin 
	 w_r = 24'b 000000000000000011111100;
	 w_i = 24'b 111111111111111111010011;
	 next_valid = 1'b1;
	 end
	11'd1054: begin 
	 w_r = 24'b 000000000000000011111100;
	 w_i = 24'b 111111111111111111010001;
	 next_valid = 1'b1;
	 end
	11'd1055: begin 
	 w_r = 24'b 000000000000000011111011;
	 w_i = 24'b 111111111111111111010000;
	 next_valid = 1'b1;
	 end
	11'd1056: begin 
	 w_r = 24'b 000000000000000011111011;
	 w_i = 24'b 111111111111111111001110;
	 next_valid = 1'b1;
	 end
	11'd1057: begin 
	 w_r = 24'b 000000000000000011111011;
	 w_i = 24'b 111111111111111111001101;
	 next_valid = 1'b1;
	 end
	11'd1058: begin 
	 w_r = 24'b 000000000000000011111010;
	 w_i = 24'b 111111111111111111001011;
	 next_valid = 1'b1;
	 end
	11'd1059: begin 
	 w_r = 24'b 000000000000000011111010;
	 w_i = 24'b 111111111111111111001001;
	 next_valid = 1'b1;
	 end
	11'd1060: begin 
	 w_r = 24'b 000000000000000011111010;
	 w_i = 24'b 111111111111111111001000;
	 next_valid = 1'b1;
	 end
	11'd1061: begin 
	 w_r = 24'b 000000000000000011111001;
	 w_i = 24'b 111111111111111111000110;
	 next_valid = 1'b1;
	 end
	11'd1062: begin 
	 w_r = 24'b 000000000000000011111001;
	 w_i = 24'b 111111111111111111000101;
	 next_valid = 1'b1;
	 end
	11'd1063: begin 
	 w_r = 24'b 000000000000000011111001;
	 w_i = 24'b 111111111111111111000011;
	 next_valid = 1'b1;
	 end
	11'd1064: begin 
	 w_r = 24'b 000000000000000011111000;
	 w_i = 24'b 111111111111111111000010;
	 next_valid = 1'b1;
	 end
	11'd1065: begin 
	 w_r = 24'b 000000000000000011111000;
	 w_i = 24'b 111111111111111111000000;
	 next_valid = 1'b1;
	 end
	11'd1066: begin 
	 w_r = 24'b 000000000000000011111000;
	 w_i = 24'b 111111111111111110111111;
	 next_valid = 1'b1;
	 end
	11'd1067: begin 
	 w_r = 24'b 000000000000000011110111;
	 w_i = 24'b 111111111111111110111101;
	 next_valid = 1'b1;
	 end
	11'd1068: begin 
	 w_r = 24'b 000000000000000011110111;
	 w_i = 24'b 111111111111111110111100;
	 next_valid = 1'b1;
	 end
	11'd1069: begin 
	 w_r = 24'b 000000000000000011110110;
	 w_i = 24'b 111111111111111110111010;
	 next_valid = 1'b1;
	 end
	11'd1070: begin 
	 w_r = 24'b 000000000000000011110110;
	 w_i = 24'b 111111111111111110111001;
	 next_valid = 1'b1;
	 end
	11'd1071: begin 
	 w_r = 24'b 000000000000000011110101;
	 w_i = 24'b 111111111111111110110111;
	 next_valid = 1'b1;
	 end
	11'd1072: begin 
	 w_r = 24'b 000000000000000011110101;
	 w_i = 24'b 111111111111111110110110;
	 next_valid = 1'b1;
	 end
	11'd1073: begin 
	 w_r = 24'b 000000000000000011110101;
	 w_i = 24'b 111111111111111110110100;
	 next_valid = 1'b1;
	 end
	11'd1074: begin 
	 w_r = 24'b 000000000000000011110100;
	 w_i = 24'b 111111111111111110110011;
	 next_valid = 1'b1;
	 end
	11'd1075: begin 
	 w_r = 24'b 000000000000000011110100;
	 w_i = 24'b 111111111111111110110001;
	 next_valid = 1'b1;
	 end
	11'd1076: begin 
	 w_r = 24'b 000000000000000011110011;
	 w_i = 24'b 111111111111111110110000;
	 next_valid = 1'b1;
	 end
	11'd1077: begin 
	 w_r = 24'b 000000000000000011110011;
	 w_i = 24'b 111111111111111110101110;
	 next_valid = 1'b1;
	 end
	11'd1078: begin 
	 w_r = 24'b 000000000000000011110010;
	 w_i = 24'b 111111111111111110101101;
	 next_valid = 1'b1;
	 end
	11'd1079: begin 
	 w_r = 24'b 000000000000000011110010;
	 w_i = 24'b 111111111111111110101011;
	 next_valid = 1'b1;
	 end
	11'd1080: begin 
	 w_r = 24'b 000000000000000011110001;
	 w_i = 24'b 111111111111111110101010;
	 next_valid = 1'b1;
	 end
	11'd1081: begin 
	 w_r = 24'b 000000000000000011110001;
	 w_i = 24'b 111111111111111110101000;
	 next_valid = 1'b1;
	 end
	11'd1082: begin 
	 w_r = 24'b 000000000000000011110000;
	 w_i = 24'b 111111111111111110100111;
	 next_valid = 1'b1;
	 end
	11'd1083: begin 
	 w_r = 24'b 000000000000000011101111;
	 w_i = 24'b 111111111111111110100101;
	 next_valid = 1'b1;
	 end
	11'd1084: begin 
	 w_r = 24'b 000000000000000011101111;
	 w_i = 24'b 111111111111111110100100;
	 next_valid = 1'b1;
	 end
	11'd1085: begin 
	 w_r = 24'b 000000000000000011101110;
	 w_i = 24'b 111111111111111110100010;
	 next_valid = 1'b1;
	 end
	11'd1086: begin 
	 w_r = 24'b 000000000000000011101110;
	 w_i = 24'b 111111111111111110100001;
	 next_valid = 1'b1;
	 end
	11'd1087: begin 
	 w_r = 24'b 000000000000000011101101;
	 w_i = 24'b 111111111111111110011111;
	 next_valid = 1'b1;
	 end
	11'd1088: begin 
	 w_r = 24'b 000000000000000011101101;
	 w_i = 24'b 111111111111111110011110;
	 next_valid = 1'b1;
	 end
	11'd1089: begin 
	 w_r = 24'b 000000000000000011101100;
	 w_i = 24'b 111111111111111110011101;
	 next_valid = 1'b1;
	 end
	11'd1090: begin 
	 w_r = 24'b 000000000000000011101011;
	 w_i = 24'b 111111111111111110011011;
	 next_valid = 1'b1;
	 end
	11'd1091: begin 
	 w_r = 24'b 000000000000000011101011;
	 w_i = 24'b 111111111111111110011010;
	 next_valid = 1'b1;
	 end
	11'd1092: begin 
	 w_r = 24'b 000000000000000011101010;
	 w_i = 24'b 111111111111111110011000;
	 next_valid = 1'b1;
	 end
	11'd1093: begin 
	 w_r = 24'b 000000000000000011101001;
	 w_i = 24'b 111111111111111110010111;
	 next_valid = 1'b1;
	 end
	11'd1094: begin 
	 w_r = 24'b 000000000000000011101001;
	 w_i = 24'b 111111111111111110010101;
	 next_valid = 1'b1;
	 end
	11'd1095: begin 
	 w_r = 24'b 000000000000000011101000;
	 w_i = 24'b 111111111111111110010100;
	 next_valid = 1'b1;
	 end
	11'd1096: begin 
	 w_r = 24'b 000000000000000011100111;
	 w_i = 24'b 111111111111111110010011;
	 next_valid = 1'b1;
	 end
	11'd1097: begin 
	 w_r = 24'b 000000000000000011100111;
	 w_i = 24'b 111111111111111110010001;
	 next_valid = 1'b1;
	 end
	11'd1098: begin 
	 w_r = 24'b 000000000000000011100110;
	 w_i = 24'b 111111111111111110010000;
	 next_valid = 1'b1;
	 end
	11'd1099: begin 
	 w_r = 24'b 000000000000000011100101;
	 w_i = 24'b 111111111111111110001110;
	 next_valid = 1'b1;
	 end
	11'd1100: begin 
	 w_r = 24'b 000000000000000011100101;
	 w_i = 24'b 111111111111111110001101;
	 next_valid = 1'b1;
	 end
	11'd1101: begin 
	 w_r = 24'b 000000000000000011100100;
	 w_i = 24'b 111111111111111110001011;
	 next_valid = 1'b1;
	 end
	11'd1102: begin 
	 w_r = 24'b 000000000000000011100011;
	 w_i = 24'b 111111111111111110001010;
	 next_valid = 1'b1;
	 end
	11'd1103: begin 
	 w_r = 24'b 000000000000000011100011;
	 w_i = 24'b 111111111111111110001001;
	 next_valid = 1'b1;
	 end
	11'd1104: begin 
	 w_r = 24'b 000000000000000011100010;
	 w_i = 24'b 111111111111111110000111;
	 next_valid = 1'b1;
	 end
	11'd1105: begin 
	 w_r = 24'b 000000000000000011100001;
	 w_i = 24'b 111111111111111110000110;
	 next_valid = 1'b1;
	 end
	11'd1106: begin 
	 w_r = 24'b 000000000000000011100000;
	 w_i = 24'b 111111111111111110000101;
	 next_valid = 1'b1;
	 end
	11'd1107: begin 
	 w_r = 24'b 000000000000000011100000;
	 w_i = 24'b 111111111111111110000011;
	 next_valid = 1'b1;
	 end
	11'd1108: begin 
	 w_r = 24'b 000000000000000011011111;
	 w_i = 24'b 111111111111111110000010;
	 next_valid = 1'b1;
	 end
	11'd1109: begin 
	 w_r = 24'b 000000000000000011011110;
	 w_i = 24'b 111111111111111110000000;
	 next_valid = 1'b1;
	 end
	11'd1110: begin 
	 w_r = 24'b 000000000000000011011101;
	 w_i = 24'b 111111111111111101111111;
	 next_valid = 1'b1;
	 end
	11'd1111: begin 
	 w_r = 24'b 000000000000000011011100;
	 w_i = 24'b 111111111111111101111110;
	 next_valid = 1'b1;
	 end
	11'd1112: begin 
	 w_r = 24'b 000000000000000011011100;
	 w_i = 24'b 111111111111111101111100;
	 next_valid = 1'b1;
	 end
	11'd1113: begin 
	 w_r = 24'b 000000000000000011011011;
	 w_i = 24'b 111111111111111101111011;
	 next_valid = 1'b1;
	 end
	11'd1114: begin 
	 w_r = 24'b 000000000000000011011010;
	 w_i = 24'b 111111111111111101111010;
	 next_valid = 1'b1;
	 end
	11'd1115: begin 
	 w_r = 24'b 000000000000000011011001;
	 w_i = 24'b 111111111111111101111000;
	 next_valid = 1'b1;
	 end
	11'd1116: begin 
	 w_r = 24'b 000000000000000011011000;
	 w_i = 24'b 111111111111111101110111;
	 next_valid = 1'b1;
	 end
	11'd1117: begin 
	 w_r = 24'b 000000000000000011010111;
	 w_i = 24'b 111111111111111101110110;
	 next_valid = 1'b1;
	 end
	11'd1118: begin 
	 w_r = 24'b 000000000000000011010111;
	 w_i = 24'b 111111111111111101110100;
	 next_valid = 1'b1;
	 end
	11'd1119: begin 
	 w_r = 24'b 000000000000000011010110;
	 w_i = 24'b 111111111111111101110011;
	 next_valid = 1'b1;
	 end
	11'd1120: begin 
	 w_r = 24'b 000000000000000011010101;
	 w_i = 24'b 111111111111111101110010;
	 next_valid = 1'b1;
	 end
	11'd1121: begin 
	 w_r = 24'b 000000000000000011010100;
	 w_i = 24'b 111111111111111101110000;
	 next_valid = 1'b1;
	 end
	11'd1122: begin 
	 w_r = 24'b 000000000000000011010011;
	 w_i = 24'b 111111111111111101101111;
	 next_valid = 1'b1;
	 end
	11'd1123: begin 
	 w_r = 24'b 000000000000000011010010;
	 w_i = 24'b 111111111111111101101110;
	 next_valid = 1'b1;
	 end
	11'd1124: begin 
	 w_r = 24'b 000000000000000011010001;
	 w_i = 24'b 111111111111111101101101;
	 next_valid = 1'b1;
	 end
	11'd1125: begin 
	 w_r = 24'b 000000000000000011010000;
	 w_i = 24'b 111111111111111101101011;
	 next_valid = 1'b1;
	 end
	11'd1126: begin 
	 w_r = 24'b 000000000000000011001111;
	 w_i = 24'b 111111111111111101101010;
	 next_valid = 1'b1;
	 end
	11'd1127: begin 
	 w_r = 24'b 000000000000000011001111;
	 w_i = 24'b 111111111111111101101001;
	 next_valid = 1'b1;
	 end
	11'd1128: begin 
	 w_r = 24'b 000000000000000011001110;
	 w_i = 24'b 111111111111111101101000;
	 next_valid = 1'b1;
	 end
	11'd1129: begin 
	 w_r = 24'b 000000000000000011001101;
	 w_i = 24'b 111111111111111101100110;
	 next_valid = 1'b1;
	 end
	11'd1130: begin 
	 w_r = 24'b 000000000000000011001100;
	 w_i = 24'b 111111111111111101100101;
	 next_valid = 1'b1;
	 end
	11'd1131: begin 
	 w_r = 24'b 000000000000000011001011;
	 w_i = 24'b 111111111111111101100100;
	 next_valid = 1'b1;
	 end
	11'd1132: begin 
	 w_r = 24'b 000000000000000011001010;
	 w_i = 24'b 111111111111111101100011;
	 next_valid = 1'b1;
	 end
	11'd1133: begin 
	 w_r = 24'b 000000000000000011001001;
	 w_i = 24'b 111111111111111101100001;
	 next_valid = 1'b1;
	 end
	11'd1134: begin 
	 w_r = 24'b 000000000000000011001000;
	 w_i = 24'b 111111111111111101100000;
	 next_valid = 1'b1;
	 end
	11'd1135: begin 
	 w_r = 24'b 000000000000000011000111;
	 w_i = 24'b 111111111111111101011111;
	 next_valid = 1'b1;
	 end
	11'd1136: begin 
	 w_r = 24'b 000000000000000011000110;
	 w_i = 24'b 111111111111111101011110;
	 next_valid = 1'b1;
	 end
	11'd1137: begin 
	 w_r = 24'b 000000000000000011000101;
	 w_i = 24'b 111111111111111101011100;
	 next_valid = 1'b1;
	 end
	11'd1138: begin 
	 w_r = 24'b 000000000000000011000100;
	 w_i = 24'b 111111111111111101011011;
	 next_valid = 1'b1;
	 end
	11'd1139: begin 
	 w_r = 24'b 000000000000000011000011;
	 w_i = 24'b 111111111111111101011010;
	 next_valid = 1'b1;
	 end
	11'd1140: begin 
	 w_r = 24'b 000000000000000011000010;
	 w_i = 24'b 111111111111111101011001;
	 next_valid = 1'b1;
	 end
	11'd1141: begin 
	 w_r = 24'b 000000000000000011000001;
	 w_i = 24'b 111111111111111101011000;
	 next_valid = 1'b1;
	 end
	11'd1142: begin 
	 w_r = 24'b 000000000000000011000000;
	 w_i = 24'b 111111111111111101010110;
	 next_valid = 1'b1;
	 end
	11'd1143: begin 
	 w_r = 24'b 000000000000000010111111;
	 w_i = 24'b 111111111111111101010101;
	 next_valid = 1'b1;
	 end
	11'd1144: begin 
	 w_r = 24'b 000000000000000010111110;
	 w_i = 24'b 111111111111111101010100;
	 next_valid = 1'b1;
	 end
	11'd1145: begin 
	 w_r = 24'b 000000000000000010111101;
	 w_i = 24'b 111111111111111101010011;
	 next_valid = 1'b1;
	 end
	11'd1146: begin 
	 w_r = 24'b 000000000000000010111100;
	 w_i = 24'b 111111111111111101010010;
	 next_valid = 1'b1;
	 end
	11'd1147: begin 
	 w_r = 24'b 000000000000000010111010;
	 w_i = 24'b 111111111111111101010001;
	 next_valid = 1'b1;
	 end
	11'd1148: begin 
	 w_r = 24'b 000000000000000010111001;
	 w_i = 24'b 111111111111111101001111;
	 next_valid = 1'b1;
	 end
	11'd1149: begin 
	 w_r = 24'b 000000000000000010111000;
	 w_i = 24'b 111111111111111101001110;
	 next_valid = 1'b1;
	 end
	11'd1150: begin 
	 w_r = 24'b 000000000000000010110111;
	 w_i = 24'b 111111111111111101001101;
	 next_valid = 1'b1;
	 end
	11'd1151: begin 
	 w_r = 24'b 000000000000000010110110;
	 w_i = 24'b 111111111111111101001100;
	 next_valid = 1'b1;
	 end
	11'd1152: begin 
	 w_r = 24'b 000000000000000010110101;
	 w_i = 24'b 111111111111111101001011;
	 next_valid = 1'b1;
	 end
	11'd1153: begin 
	 w_r = 24'b 000000000000000010110100;
	 w_i = 24'b 111111111111111101001010;
	 next_valid = 1'b1;
	 end
	11'd1154: begin 
	 w_r = 24'b 000000000000000010110011;
	 w_i = 24'b 111111111111111101001001;
	 next_valid = 1'b1;
	 end
	11'd1155: begin 
	 w_r = 24'b 000000000000000010110010;
	 w_i = 24'b 111111111111111101001000;
	 next_valid = 1'b1;
	 end
	11'd1156: begin 
	 w_r = 24'b 000000000000000010110001;
	 w_i = 24'b 111111111111111101000111;
	 next_valid = 1'b1;
	 end
	11'd1157: begin 
	 w_r = 24'b 000000000000000010101111;
	 w_i = 24'b 111111111111111101000110;
	 next_valid = 1'b1;
	 end
	11'd1158: begin 
	 w_r = 24'b 000000000000000010101110;
	 w_i = 24'b 111111111111111101000100;
	 next_valid = 1'b1;
	 end
	11'd1159: begin 
	 w_r = 24'b 000000000000000010101101;
	 w_i = 24'b 111111111111111101000011;
	 next_valid = 1'b1;
	 end
	11'd1160: begin 
	 w_r = 24'b 000000000000000010101100;
	 w_i = 24'b 111111111111111101000010;
	 next_valid = 1'b1;
	 end
	11'd1161: begin 
	 w_r = 24'b 000000000000000010101011;
	 w_i = 24'b 111111111111111101000001;
	 next_valid = 1'b1;
	 end
	11'd1162: begin 
	 w_r = 24'b 000000000000000010101010;
	 w_i = 24'b 111111111111111101000000;
	 next_valid = 1'b1;
	 end
	11'd1163: begin 
	 w_r = 24'b 000000000000000010101000;
	 w_i = 24'b 111111111111111100111111;
	 next_valid = 1'b1;
	 end
	11'd1164: begin 
	 w_r = 24'b 000000000000000010100111;
	 w_i = 24'b 111111111111111100111110;
	 next_valid = 1'b1;
	 end
	11'd1165: begin 
	 w_r = 24'b 000000000000000010100110;
	 w_i = 24'b 111111111111111100111101;
	 next_valid = 1'b1;
	 end
	11'd1166: begin 
	 w_r = 24'b 000000000000000010100101;
	 w_i = 24'b 111111111111111100111100;
	 next_valid = 1'b1;
	 end
	11'd1167: begin 
	 w_r = 24'b 000000000000000010100100;
	 w_i = 24'b 111111111111111100111011;
	 next_valid = 1'b1;
	 end
	11'd1168: begin 
	 w_r = 24'b 000000000000000010100010;
	 w_i = 24'b 111111111111111100111010;
	 next_valid = 1'b1;
	 end
	11'd1169: begin 
	 w_r = 24'b 000000000000000010100001;
	 w_i = 24'b 111111111111111100111001;
	 next_valid = 1'b1;
	 end
	11'd1170: begin 
	 w_r = 24'b 000000000000000010100000;
	 w_i = 24'b 111111111111111100111000;
	 next_valid = 1'b1;
	 end
	11'd1171: begin 
	 w_r = 24'b 000000000000000010011111;
	 w_i = 24'b 111111111111111100110111;
	 next_valid = 1'b1;
	 end
	11'd1172: begin 
	 w_r = 24'b 000000000000000010011101;
	 w_i = 24'b 111111111111111100110110;
	 next_valid = 1'b1;
	 end
	11'd1173: begin 
	 w_r = 24'b 000000000000000010011100;
	 w_i = 24'b 111111111111111100110101;
	 next_valid = 1'b1;
	 end
	11'd1174: begin 
	 w_r = 24'b 000000000000000010011011;
	 w_i = 24'b 111111111111111100110100;
	 next_valid = 1'b1;
	 end
	11'd1175: begin 
	 w_r = 24'b 000000000000000010011010;
	 w_i = 24'b 111111111111111100110011;
	 next_valid = 1'b1;
	 end
	11'd1176: begin 
	 w_r = 24'b 000000000000000010011000;
	 w_i = 24'b 111111111111111100110010;
	 next_valid = 1'b1;
	 end
	11'd1177: begin 
	 w_r = 24'b 000000000000000010010111;
	 w_i = 24'b 111111111111111100110001;
	 next_valid = 1'b1;
	 end
	11'd1178: begin 
	 w_r = 24'b 000000000000000010010110;
	 w_i = 24'b 111111111111111100110001;
	 next_valid = 1'b1;
	 end
	11'd1179: begin 
	 w_r = 24'b 000000000000000010010101;
	 w_i = 24'b 111111111111111100110000;
	 next_valid = 1'b1;
	 end
	11'd1180: begin 
	 w_r = 24'b 000000000000000010010011;
	 w_i = 24'b 111111111111111100101111;
	 next_valid = 1'b1;
	 end
	11'd1181: begin 
	 w_r = 24'b 000000000000000010010010;
	 w_i = 24'b 111111111111111100101110;
	 next_valid = 1'b1;
	 end
	11'd1182: begin 
	 w_r = 24'b 000000000000000010010001;
	 w_i = 24'b 111111111111111100101101;
	 next_valid = 1'b1;
	 end
	11'd1183: begin 
	 w_r = 24'b 000000000000000010010000;
	 w_i = 24'b 111111111111111100101100;
	 next_valid = 1'b1;
	 end
	11'd1184: begin 
	 w_r = 24'b 000000000000000010001110;
	 w_i = 24'b 111111111111111100101011;
	 next_valid = 1'b1;
	 end
	11'd1185: begin 
	 w_r = 24'b 000000000000000010001101;
	 w_i = 24'b 111111111111111100101010;
	 next_valid = 1'b1;
	 end
	11'd1186: begin 
	 w_r = 24'b 000000000000000010001100;
	 w_i = 24'b 111111111111111100101001;
	 next_valid = 1'b1;
	 end
	11'd1187: begin 
	 w_r = 24'b 000000000000000010001010;
	 w_i = 24'b 111111111111111100101001;
	 next_valid = 1'b1;
	 end
	11'd1188: begin 
	 w_r = 24'b 000000000000000010001001;
	 w_i = 24'b 111111111111111100101000;
	 next_valid = 1'b1;
	 end
	11'd1189: begin 
	 w_r = 24'b 000000000000000010001000;
	 w_i = 24'b 111111111111111100100111;
	 next_valid = 1'b1;
	 end
	11'd1190: begin 
	 w_r = 24'b 000000000000000010000110;
	 w_i = 24'b 111111111111111100100110;
	 next_valid = 1'b1;
	 end
	11'd1191: begin 
	 w_r = 24'b 000000000000000010000101;
	 w_i = 24'b 111111111111111100100101;
	 next_valid = 1'b1;
	 end
	11'd1192: begin 
	 w_r = 24'b 000000000000000010000100;
	 w_i = 24'b 111111111111111100100100;
	 next_valid = 1'b1;
	 end
	11'd1193: begin 
	 w_r = 24'b 000000000000000010000010;
	 w_i = 24'b 111111111111111100100100;
	 next_valid = 1'b1;
	 end
	11'd1194: begin 
	 w_r = 24'b 000000000000000010000001;
	 w_i = 24'b 111111111111111100100011;
	 next_valid = 1'b1;
	 end
	11'd1195: begin 
	 w_r = 24'b 000000000000000010000000;
	 w_i = 24'b 111111111111111100100010;
	 next_valid = 1'b1;
	 end
	11'd1196: begin 
	 w_r = 24'b 000000000000000001111110;
	 w_i = 24'b 111111111111111100100001;
	 next_valid = 1'b1;
	 end
	11'd1197: begin 
	 w_r = 24'b 000000000000000001111101;
	 w_i = 24'b 111111111111111100100000;
	 next_valid = 1'b1;
	 end
	11'd1198: begin 
	 w_r = 24'b 000000000000000001111011;
	 w_i = 24'b 111111111111111100100000;
	 next_valid = 1'b1;
	 end
	11'd1199: begin 
	 w_r = 24'b 000000000000000001111010;
	 w_i = 24'b 111111111111111100011111;
	 next_valid = 1'b1;
	 end
	11'd1200: begin 
	 w_r = 24'b 000000000000000001111001;
	 w_i = 24'b 111111111111111100011110;
	 next_valid = 1'b1;
	 end
	11'd1201: begin 
	 w_r = 24'b 000000000000000001110111;
	 w_i = 24'b 111111111111111100011101;
	 next_valid = 1'b1;
	 end
	11'd1202: begin 
	 w_r = 24'b 000000000000000001110110;
	 w_i = 24'b 111111111111111100011101;
	 next_valid = 1'b1;
	 end
	11'd1203: begin 
	 w_r = 24'b 000000000000000001110101;
	 w_i = 24'b 111111111111111100011100;
	 next_valid = 1'b1;
	 end
	11'd1204: begin 
	 w_r = 24'b 000000000000000001110011;
	 w_i = 24'b 111111111111111100011011;
	 next_valid = 1'b1;
	 end
	11'd1205: begin 
	 w_r = 24'b 000000000000000001110010;
	 w_i = 24'b 111111111111111100011011;
	 next_valid = 1'b1;
	 end
	11'd1206: begin 
	 w_r = 24'b 000000000000000001110000;
	 w_i = 24'b 111111111111111100011010;
	 next_valid = 1'b1;
	 end
	11'd1207: begin 
	 w_r = 24'b 000000000000000001101111;
	 w_i = 24'b 111111111111111100011001;
	 next_valid = 1'b1;
	 end
	11'd1208: begin 
	 w_r = 24'b 000000000000000001101101;
	 w_i = 24'b 111111111111111100011001;
	 next_valid = 1'b1;
	 end
	11'd1209: begin 
	 w_r = 24'b 000000000000000001101100;
	 w_i = 24'b 111111111111111100011000;
	 next_valid = 1'b1;
	 end
	11'd1210: begin 
	 w_r = 24'b 000000000000000001101011;
	 w_i = 24'b 111111111111111100010111;
	 next_valid = 1'b1;
	 end
	11'd1211: begin 
	 w_r = 24'b 000000000000000001101001;
	 w_i = 24'b 111111111111111100010111;
	 next_valid = 1'b1;
	 end
	11'd1212: begin 
	 w_r = 24'b 000000000000000001101000;
	 w_i = 24'b 111111111111111100010110;
	 next_valid = 1'b1;
	 end
	11'd1213: begin 
	 w_r = 24'b 000000000000000001100110;
	 w_i = 24'b 111111111111111100010101;
	 next_valid = 1'b1;
	 end
	11'd1214: begin 
	 w_r = 24'b 000000000000000001100101;
	 w_i = 24'b 111111111111111100010101;
	 next_valid = 1'b1;
	 end
	11'd1215: begin 
	 w_r = 24'b 000000000000000001100011;
	 w_i = 24'b 111111111111111100010100;
	 next_valid = 1'b1;
	 end
	11'd1216: begin 
	 w_r = 24'b 000000000000000001100010;
	 w_i = 24'b 111111111111111100010011;
	 next_valid = 1'b1;
	 end
	11'd1217: begin 
	 w_r = 24'b 000000000000000001100001;
	 w_i = 24'b 111111111111111100010011;
	 next_valid = 1'b1;
	 end
	11'd1218: begin 
	 w_r = 24'b 000000000000000001011111;
	 w_i = 24'b 111111111111111100010010;
	 next_valid = 1'b1;
	 end
	11'd1219: begin 
	 w_r = 24'b 000000000000000001011110;
	 w_i = 24'b 111111111111111100010010;
	 next_valid = 1'b1;
	 end
	11'd1220: begin 
	 w_r = 24'b 000000000000000001011100;
	 w_i = 24'b 111111111111111100010001;
	 next_valid = 1'b1;
	 end
	11'd1221: begin 
	 w_r = 24'b 000000000000000001011011;
	 w_i = 24'b 111111111111111100010001;
	 next_valid = 1'b1;
	 end
	11'd1222: begin 
	 w_r = 24'b 000000000000000001011001;
	 w_i = 24'b 111111111111111100010000;
	 next_valid = 1'b1;
	 end
	11'd1223: begin 
	 w_r = 24'b 000000000000000001011000;
	 w_i = 24'b 111111111111111100001111;
	 next_valid = 1'b1;
	 end
	11'd1224: begin 
	 w_r = 24'b 000000000000000001010110;
	 w_i = 24'b 111111111111111100001111;
	 next_valid = 1'b1;
	 end
	11'd1225: begin 
	 w_r = 24'b 000000000000000001010101;
	 w_i = 24'b 111111111111111100001110;
	 next_valid = 1'b1;
	 end
	11'd1226: begin 
	 w_r = 24'b 000000000000000001010011;
	 w_i = 24'b 111111111111111100001110;
	 next_valid = 1'b1;
	 end
	11'd1227: begin 
	 w_r = 24'b 000000000000000001010010;
	 w_i = 24'b 111111111111111100001101;
	 next_valid = 1'b1;
	 end
	11'd1228: begin 
	 w_r = 24'b 000000000000000001010000;
	 w_i = 24'b 111111111111111100001101;
	 next_valid = 1'b1;
	 end
	11'd1229: begin 
	 w_r = 24'b 000000000000000001001111;
	 w_i = 24'b 111111111111111100001100;
	 next_valid = 1'b1;
	 end
	11'd1230: begin 
	 w_r = 24'b 000000000000000001001101;
	 w_i = 24'b 111111111111111100001100;
	 next_valid = 1'b1;
	 end
	11'd1231: begin 
	 w_r = 24'b 000000000000000001001100;
	 w_i = 24'b 111111111111111100001011;
	 next_valid = 1'b1;
	 end
	11'd1232: begin 
	 w_r = 24'b 000000000000000001001010;
	 w_i = 24'b 111111111111111100001011;
	 next_valid = 1'b1;
	 end
	11'd1233: begin 
	 w_r = 24'b 000000000000000001001001;
	 w_i = 24'b 111111111111111100001011;
	 next_valid = 1'b1;
	 end
	11'd1234: begin 
	 w_r = 24'b 000000000000000001000111;
	 w_i = 24'b 111111111111111100001010;
	 next_valid = 1'b1;
	 end
	11'd1235: begin 
	 w_r = 24'b 000000000000000001000110;
	 w_i = 24'b 111111111111111100001010;
	 next_valid = 1'b1;
	 end
	11'd1236: begin 
	 w_r = 24'b 000000000000000001000100;
	 w_i = 24'b 111111111111111100001001;
	 next_valid = 1'b1;
	 end
	11'd1237: begin 
	 w_r = 24'b 000000000000000001000011;
	 w_i = 24'b 111111111111111100001001;
	 next_valid = 1'b1;
	 end
	11'd1238: begin 
	 w_r = 24'b 000000000000000001000001;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	11'd1239: begin 
	 w_r = 24'b 000000000000000001000000;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	11'd1240: begin 
	 w_r = 24'b 000000000000000000111110;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	11'd1241: begin 
	 w_r = 24'b 000000000000000000111101;
	 w_i = 24'b 111111111111111100000111;
	 next_valid = 1'b1;
	 end
	11'd1242: begin 
	 w_r = 24'b 000000000000000000111011;
	 w_i = 24'b 111111111111111100000111;
	 next_valid = 1'b1;
	 end
	11'd1243: begin 
	 w_r = 24'b 000000000000000000111010;
	 w_i = 24'b 111111111111111100000111;
	 next_valid = 1'b1;
	 end
	11'd1244: begin 
	 w_r = 24'b 000000000000000000111000;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	11'd1245: begin 
	 w_r = 24'b 000000000000000000110111;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	11'd1246: begin 
	 w_r = 24'b 000000000000000000110101;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	11'd1247: begin 
	 w_r = 24'b 000000000000000000110011;
	 w_i = 24'b 111111111111111100000101;
	 next_valid = 1'b1;
	 end
	11'd1248: begin 
	 w_r = 24'b 000000000000000000110010;
	 w_i = 24'b 111111111111111100000101;
	 next_valid = 1'b1;
	 end
	11'd1249: begin 
	 w_r = 24'b 000000000000000000110000;
	 w_i = 24'b 111111111111111100000101;
	 next_valid = 1'b1;
	 end
	11'd1250: begin 
	 w_r = 24'b 000000000000000000101111;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	11'd1251: begin 
	 w_r = 24'b 000000000000000000101101;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	11'd1252: begin 
	 w_r = 24'b 000000000000000000101100;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	11'd1253: begin 
	 w_r = 24'b 000000000000000000101010;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	11'd1254: begin 
	 w_r = 24'b 000000000000000000101001;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	11'd1255: begin 
	 w_r = 24'b 000000000000000000100111;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	11'd1256: begin 
	 w_r = 24'b 000000000000000000100110;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	11'd1257: begin 
	 w_r = 24'b 000000000000000000100100;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	11'd1258: begin 
	 w_r = 24'b 000000000000000000100010;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	11'd1259: begin 
	 w_r = 24'b 000000000000000000100001;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	11'd1260: begin 
	 w_r = 24'b 000000000000000000011111;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	11'd1261: begin 
	 w_r = 24'b 000000000000000000011110;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	11'd1262: begin 
	 w_r = 24'b 000000000000000000011100;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	11'd1263: begin 
	 w_r = 24'b 000000000000000000011011;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1264: begin 
	 w_r = 24'b 000000000000000000011001;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1265: begin 
	 w_r = 24'b 000000000000000000011000;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1266: begin 
	 w_r = 24'b 000000000000000000010110;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1267: begin 
	 w_r = 24'b 000000000000000000010100;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1268: begin 
	 w_r = 24'b 000000000000000000010011;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1269: begin 
	 w_r = 24'b 000000000000000000010001;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1270: begin 
	 w_r = 24'b 000000000000000000010000;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1271: begin 
	 w_r = 24'b 000000000000000000001110;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1272: begin 
	 w_r = 24'b 000000000000000000001101;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1273: begin 
	 w_r = 24'b 000000000000000000001011;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1274: begin 
	 w_r = 24'b 000000000000000000001001;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1275: begin 
	 w_r = 24'b 000000000000000000001000;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1276: begin 
	 w_r = 24'b 000000000000000000000110;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1277: begin 
	 w_r = 24'b 000000000000000000000101;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1278: begin 
	 w_r = 24'b 000000000000000000000011;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1279: begin 
	 w_r = 24'b 000000000000000000000010;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1280: begin 
	 w_r = 24'b 000000000000000000000000;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1281: begin 
	 w_r = 24'b 111111111111111111111110;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1282: begin 
	 w_r = 24'b 111111111111111111111101;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1283: begin 
	 w_r = 24'b 111111111111111111111011;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1284: begin 
	 w_r = 24'b 111111111111111111111010;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1285: begin 
	 w_r = 24'b 111111111111111111111000;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1286: begin 
	 w_r = 24'b 111111111111111111110111;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1287: begin 
	 w_r = 24'b 111111111111111111110101;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1288: begin 
	 w_r = 24'b 111111111111111111110011;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1289: begin 
	 w_r = 24'b 111111111111111111110010;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1290: begin 
	 w_r = 24'b 111111111111111111110000;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	11'd1291: begin 
	 w_r = 24'b 111111111111111111101111;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1292: begin 
	 w_r = 24'b 111111111111111111101101;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1293: begin 
	 w_r = 24'b 111111111111111111101100;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1294: begin 
	 w_r = 24'b 111111111111111111101010;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1295: begin 
	 w_r = 24'b 111111111111111111101000;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1296: begin 
	 w_r = 24'b 111111111111111111100111;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1297: begin 
	 w_r = 24'b 111111111111111111100101;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	11'd1298: begin 
	 w_r = 24'b 111111111111111111100100;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	11'd1299: begin 
	 w_r = 24'b 111111111111111111100010;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	11'd1300: begin 
	 w_r = 24'b 111111111111111111100001;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	11'd1301: begin 
	 w_r = 24'b 111111111111111111011111;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	11'd1302: begin 
	 w_r = 24'b 111111111111111111011110;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	11'd1303: begin 
	 w_r = 24'b 111111111111111111011100;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	11'd1304: begin 
	 w_r = 24'b 111111111111111111011010;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	11'd1305: begin 
	 w_r = 24'b 111111111111111111011001;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	11'd1306: begin 
	 w_r = 24'b 111111111111111111010111;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	11'd1307: begin 
	 w_r = 24'b 111111111111111111010110;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	11'd1308: begin 
	 w_r = 24'b 111111111111111111010100;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	11'd1309: begin 
	 w_r = 24'b 111111111111111111010011;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	11'd1310: begin 
	 w_r = 24'b 111111111111111111010001;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	11'd1311: begin 
	 w_r = 24'b 111111111111111111010000;
	 w_i = 24'b 111111111111111100000101;
	 next_valid = 1'b1;
	 end
	11'd1312: begin 
	 w_r = 24'b 111111111111111111001110;
	 w_i = 24'b 111111111111111100000101;
	 next_valid = 1'b1;
	 end
	11'd1313: begin 
	 w_r = 24'b 111111111111111111001101;
	 w_i = 24'b 111111111111111100000101;
	 next_valid = 1'b1;
	 end
	11'd1314: begin 
	 w_r = 24'b 111111111111111111001011;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	11'd1315: begin 
	 w_r = 24'b 111111111111111111001001;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	11'd1316: begin 
	 w_r = 24'b 111111111111111111001000;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	11'd1317: begin 
	 w_r = 24'b 111111111111111111000110;
	 w_i = 24'b 111111111111111100000111;
	 next_valid = 1'b1;
	 end
	11'd1318: begin 
	 w_r = 24'b 111111111111111111000101;
	 w_i = 24'b 111111111111111100000111;
	 next_valid = 1'b1;
	 end
	11'd1319: begin 
	 w_r = 24'b 111111111111111111000011;
	 w_i = 24'b 111111111111111100000111;
	 next_valid = 1'b1;
	 end
	11'd1320: begin 
	 w_r = 24'b 111111111111111111000010;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	11'd1321: begin 
	 w_r = 24'b 111111111111111111000000;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	11'd1322: begin 
	 w_r = 24'b 111111111111111110111111;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	11'd1323: begin 
	 w_r = 24'b 111111111111111110111101;
	 w_i = 24'b 111111111111111100001001;
	 next_valid = 1'b1;
	 end
	11'd1324: begin 
	 w_r = 24'b 111111111111111110111100;
	 w_i = 24'b 111111111111111100001001;
	 next_valid = 1'b1;
	 end
	11'd1325: begin 
	 w_r = 24'b 111111111111111110111010;
	 w_i = 24'b 111111111111111100001010;
	 next_valid = 1'b1;
	 end
	11'd1326: begin 
	 w_r = 24'b 111111111111111110111001;
	 w_i = 24'b 111111111111111100001010;
	 next_valid = 1'b1;
	 end
	11'd1327: begin 
	 w_r = 24'b 111111111111111110110111;
	 w_i = 24'b 111111111111111100001011;
	 next_valid = 1'b1;
	 end
	11'd1328: begin 
	 w_r = 24'b 111111111111111110110110;
	 w_i = 24'b 111111111111111100001011;
	 next_valid = 1'b1;
	 end
	11'd1329: begin 
	 w_r = 24'b 111111111111111110110100;
	 w_i = 24'b 111111111111111100001011;
	 next_valid = 1'b1;
	 end
	11'd1330: begin 
	 w_r = 24'b 111111111111111110110011;
	 w_i = 24'b 111111111111111100001100;
	 next_valid = 1'b1;
	 end
	11'd1331: begin 
	 w_r = 24'b 111111111111111110110001;
	 w_i = 24'b 111111111111111100001100;
	 next_valid = 1'b1;
	 end
	11'd1332: begin 
	 w_r = 24'b 111111111111111110110000;
	 w_i = 24'b 111111111111111100001101;
	 next_valid = 1'b1;
	 end
	11'd1333: begin 
	 w_r = 24'b 111111111111111110101110;
	 w_i = 24'b 111111111111111100001101;
	 next_valid = 1'b1;
	 end
	11'd1334: begin 
	 w_r = 24'b 111111111111111110101101;
	 w_i = 24'b 111111111111111100001110;
	 next_valid = 1'b1;
	 end
	11'd1335: begin 
	 w_r = 24'b 111111111111111110101011;
	 w_i = 24'b 111111111111111100001110;
	 next_valid = 1'b1;
	 end
	11'd1336: begin 
	 w_r = 24'b 111111111111111110101010;
	 w_i = 24'b 111111111111111100001111;
	 next_valid = 1'b1;
	 end
	11'd1337: begin 
	 w_r = 24'b 111111111111111110101000;
	 w_i = 24'b 111111111111111100001111;
	 next_valid = 1'b1;
	 end
	11'd1338: begin 
	 w_r = 24'b 111111111111111110100111;
	 w_i = 24'b 111111111111111100010000;
	 next_valid = 1'b1;
	 end
	11'd1339: begin 
	 w_r = 24'b 111111111111111110100101;
	 w_i = 24'b 111111111111111100010001;
	 next_valid = 1'b1;
	 end
	11'd1340: begin 
	 w_r = 24'b 111111111111111110100100;
	 w_i = 24'b 111111111111111100010001;
	 next_valid = 1'b1;
	 end
	11'd1341: begin 
	 w_r = 24'b 111111111111111110100010;
	 w_i = 24'b 111111111111111100010010;
	 next_valid = 1'b1;
	 end
	11'd1342: begin 
	 w_r = 24'b 111111111111111110100001;
	 w_i = 24'b 111111111111111100010010;
	 next_valid = 1'b1;
	 end
	11'd1343: begin 
	 w_r = 24'b 111111111111111110011111;
	 w_i = 24'b 111111111111111100010011;
	 next_valid = 1'b1;
	 end
	11'd1344: begin 
	 w_r = 24'b 111111111111111110011110;
	 w_i = 24'b 111111111111111100010011;
	 next_valid = 1'b1;
	 end
	11'd1345: begin 
	 w_r = 24'b 111111111111111110011101;
	 w_i = 24'b 111111111111111100010100;
	 next_valid = 1'b1;
	 end
	11'd1346: begin 
	 w_r = 24'b 111111111111111110011011;
	 w_i = 24'b 111111111111111100010101;
	 next_valid = 1'b1;
	 end
	11'd1347: begin 
	 w_r = 24'b 111111111111111110011010;
	 w_i = 24'b 111111111111111100010101;
	 next_valid = 1'b1;
	 end
	11'd1348: begin 
	 w_r = 24'b 111111111111111110011000;
	 w_i = 24'b 111111111111111100010110;
	 next_valid = 1'b1;
	 end
	11'd1349: begin 
	 w_r = 24'b 111111111111111110010111;
	 w_i = 24'b 111111111111111100010111;
	 next_valid = 1'b1;
	 end
	11'd1350: begin 
	 w_r = 24'b 111111111111111110010101;
	 w_i = 24'b 111111111111111100010111;
	 next_valid = 1'b1;
	 end
	11'd1351: begin 
	 w_r = 24'b 111111111111111110010100;
	 w_i = 24'b 111111111111111100011000;
	 next_valid = 1'b1;
	 end
	11'd1352: begin 
	 w_r = 24'b 111111111111111110010011;
	 w_i = 24'b 111111111111111100011001;
	 next_valid = 1'b1;
	 end
	11'd1353: begin 
	 w_r = 24'b 111111111111111110010001;
	 w_i = 24'b 111111111111111100011001;
	 next_valid = 1'b1;
	 end
	11'd1354: begin 
	 w_r = 24'b 111111111111111110010000;
	 w_i = 24'b 111111111111111100011010;
	 next_valid = 1'b1;
	 end
	11'd1355: begin 
	 w_r = 24'b 111111111111111110001110;
	 w_i = 24'b 111111111111111100011011;
	 next_valid = 1'b1;
	 end
	11'd1356: begin 
	 w_r = 24'b 111111111111111110001101;
	 w_i = 24'b 111111111111111100011011;
	 next_valid = 1'b1;
	 end
	11'd1357: begin 
	 w_r = 24'b 111111111111111110001011;
	 w_i = 24'b 111111111111111100011100;
	 next_valid = 1'b1;
	 end
	11'd1358: begin 
	 w_r = 24'b 111111111111111110001010;
	 w_i = 24'b 111111111111111100011101;
	 next_valid = 1'b1;
	 end
	11'd1359: begin 
	 w_r = 24'b 111111111111111110001001;
	 w_i = 24'b 111111111111111100011101;
	 next_valid = 1'b1;
	 end
	11'd1360: begin 
	 w_r = 24'b 111111111111111110000111;
	 w_i = 24'b 111111111111111100011110;
	 next_valid = 1'b1;
	 end
	11'd1361: begin 
	 w_r = 24'b 111111111111111110000110;
	 w_i = 24'b 111111111111111100011111;
	 next_valid = 1'b1;
	 end
	11'd1362: begin 
	 w_r = 24'b 111111111111111110000101;
	 w_i = 24'b 111111111111111100100000;
	 next_valid = 1'b1;
	 end
	11'd1363: begin 
	 w_r = 24'b 111111111111111110000011;
	 w_i = 24'b 111111111111111100100000;
	 next_valid = 1'b1;
	 end
	11'd1364: begin 
	 w_r = 24'b 111111111111111110000010;
	 w_i = 24'b 111111111111111100100001;
	 next_valid = 1'b1;
	 end
	11'd1365: begin 
	 w_r = 24'b 111111111111111110000000;
	 w_i = 24'b 111111111111111100100010;
	 next_valid = 1'b1;
	 end
	11'd1366: begin 
	 w_r = 24'b 111111111111111101111111;
	 w_i = 24'b 111111111111111100100011;
	 next_valid = 1'b1;
	 end
	11'd1367: begin 
	 w_r = 24'b 111111111111111101111110;
	 w_i = 24'b 111111111111111100100100;
	 next_valid = 1'b1;
	 end
	11'd1368: begin 
	 w_r = 24'b 111111111111111101111100;
	 w_i = 24'b 111111111111111100100100;
	 next_valid = 1'b1;
	 end
	11'd1369: begin 
	 w_r = 24'b 111111111111111101111011;
	 w_i = 24'b 111111111111111100100101;
	 next_valid = 1'b1;
	 end
	11'd1370: begin 
	 w_r = 24'b 111111111111111101111010;
	 w_i = 24'b 111111111111111100100110;
	 next_valid = 1'b1;
	 end
	11'd1371: begin 
	 w_r = 24'b 111111111111111101111000;
	 w_i = 24'b 111111111111111100100111;
	 next_valid = 1'b1;
	 end
	11'd1372: begin 
	 w_r = 24'b 111111111111111101110111;
	 w_i = 24'b 111111111111111100101000;
	 next_valid = 1'b1;
	 end
	11'd1373: begin 
	 w_r = 24'b 111111111111111101110110;
	 w_i = 24'b 111111111111111100101001;
	 next_valid = 1'b1;
	 end
	11'd1374: begin 
	 w_r = 24'b 111111111111111101110100;
	 w_i = 24'b 111111111111111100101001;
	 next_valid = 1'b1;
	 end
	11'd1375: begin 
	 w_r = 24'b 111111111111111101110011;
	 w_i = 24'b 111111111111111100101010;
	 next_valid = 1'b1;
	 end
	11'd1376: begin 
	 w_r = 24'b 111111111111111101110010;
	 w_i = 24'b 111111111111111100101011;
	 next_valid = 1'b1;
	 end
	11'd1377: begin 
	 w_r = 24'b 111111111111111101110000;
	 w_i = 24'b 111111111111111100101100;
	 next_valid = 1'b1;
	 end
	11'd1378: begin 
	 w_r = 24'b 111111111111111101101111;
	 w_i = 24'b 111111111111111100101101;
	 next_valid = 1'b1;
	 end
	11'd1379: begin 
	 w_r = 24'b 111111111111111101101110;
	 w_i = 24'b 111111111111111100101110;
	 next_valid = 1'b1;
	 end
	11'd1380: begin 
	 w_r = 24'b 111111111111111101101101;
	 w_i = 24'b 111111111111111100101111;
	 next_valid = 1'b1;
	 end
	11'd1381: begin 
	 w_r = 24'b 111111111111111101101011;
	 w_i = 24'b 111111111111111100110000;
	 next_valid = 1'b1;
	 end
	11'd1382: begin 
	 w_r = 24'b 111111111111111101101010;
	 w_i = 24'b 111111111111111100110001;
	 next_valid = 1'b1;
	 end
	11'd1383: begin 
	 w_r = 24'b 111111111111111101101001;
	 w_i = 24'b 111111111111111100110001;
	 next_valid = 1'b1;
	 end
	11'd1384: begin 
	 w_r = 24'b 111111111111111101101000;
	 w_i = 24'b 111111111111111100110010;
	 next_valid = 1'b1;
	 end
	11'd1385: begin 
	 w_r = 24'b 111111111111111101100110;
	 w_i = 24'b 111111111111111100110011;
	 next_valid = 1'b1;
	 end
	11'd1386: begin 
	 w_r = 24'b 111111111111111101100101;
	 w_i = 24'b 111111111111111100110100;
	 next_valid = 1'b1;
	 end
	11'd1387: begin 
	 w_r = 24'b 111111111111111101100100;
	 w_i = 24'b 111111111111111100110101;
	 next_valid = 1'b1;
	 end
	11'd1388: begin 
	 w_r = 24'b 111111111111111101100011;
	 w_i = 24'b 111111111111111100110110;
	 next_valid = 1'b1;
	 end
	11'd1389: begin 
	 w_r = 24'b 111111111111111101100001;
	 w_i = 24'b 111111111111111100110111;
	 next_valid = 1'b1;
	 end
	11'd1390: begin 
	 w_r = 24'b 111111111111111101100000;
	 w_i = 24'b 111111111111111100111000;
	 next_valid = 1'b1;
	 end
	11'd1391: begin 
	 w_r = 24'b 111111111111111101011111;
	 w_i = 24'b 111111111111111100111001;
	 next_valid = 1'b1;
	 end
	11'd1392: begin 
	 w_r = 24'b 111111111111111101011110;
	 w_i = 24'b 111111111111111100111010;
	 next_valid = 1'b1;
	 end
	11'd1393: begin 
	 w_r = 24'b 111111111111111101011100;
	 w_i = 24'b 111111111111111100111011;
	 next_valid = 1'b1;
	 end
	11'd1394: begin 
	 w_r = 24'b 111111111111111101011011;
	 w_i = 24'b 111111111111111100111100;
	 next_valid = 1'b1;
	 end
	11'd1395: begin 
	 w_r = 24'b 111111111111111101011010;
	 w_i = 24'b 111111111111111100111101;
	 next_valid = 1'b1;
	 end
	11'd1396: begin 
	 w_r = 24'b 111111111111111101011001;
	 w_i = 24'b 111111111111111100111110;
	 next_valid = 1'b1;
	 end
	11'd1397: begin 
	 w_r = 24'b 111111111111111101011000;
	 w_i = 24'b 111111111111111100111111;
	 next_valid = 1'b1;
	 end
	11'd1398: begin 
	 w_r = 24'b 111111111111111101010110;
	 w_i = 24'b 111111111111111101000000;
	 next_valid = 1'b1;
	 end
	11'd1399: begin 
	 w_r = 24'b 111111111111111101010101;
	 w_i = 24'b 111111111111111101000001;
	 next_valid = 1'b1;
	 end
	11'd1400: begin 
	 w_r = 24'b 111111111111111101010100;
	 w_i = 24'b 111111111111111101000010;
	 next_valid = 1'b1;
	 end
	11'd1401: begin 
	 w_r = 24'b 111111111111111101010011;
	 w_i = 24'b 111111111111111101000011;
	 next_valid = 1'b1;
	 end
	11'd1402: begin 
	 w_r = 24'b 111111111111111101010010;
	 w_i = 24'b 111111111111111101000100;
	 next_valid = 1'b1;
	 end
	11'd1403: begin 
	 w_r = 24'b 111111111111111101010001;
	 w_i = 24'b 111111111111111101000110;
	 next_valid = 1'b1;
	 end
	11'd1404: begin 
	 w_r = 24'b 111111111111111101001111;
	 w_i = 24'b 111111111111111101000111;
	 next_valid = 1'b1;
	 end
	11'd1405: begin 
	 w_r = 24'b 111111111111111101001110;
	 w_i = 24'b 111111111111111101001000;
	 next_valid = 1'b1;
	 end
	11'd1406: begin 
	 w_r = 24'b 111111111111111101001101;
	 w_i = 24'b 111111111111111101001001;
	 next_valid = 1'b1;
	 end
	11'd1407: begin 
	 w_r = 24'b 111111111111111101001100;
	 w_i = 24'b 111111111111111101001010;
	 next_valid = 1'b1;
	 end
	11'd1408: begin 
	 w_r = 24'b 111111111111111101001011;
	 w_i = 24'b 111111111111111101001011;
	 next_valid = 1'b1;
	 end
	11'd1409: begin 
	 w_r = 24'b 111111111111111101001010;
	 w_i = 24'b 111111111111111101001100;
	 next_valid = 1'b1;
	 end
	11'd1410: begin 
	 w_r = 24'b 111111111111111101001001;
	 w_i = 24'b 111111111111111101001101;
	 next_valid = 1'b1;
	 end
	11'd1411: begin 
	 w_r = 24'b 111111111111111101001000;
	 w_i = 24'b 111111111111111101001110;
	 next_valid = 1'b1;
	 end
	11'd1412: begin 
	 w_r = 24'b 111111111111111101000111;
	 w_i = 24'b 111111111111111101001111;
	 next_valid = 1'b1;
	 end
	11'd1413: begin 
	 w_r = 24'b 111111111111111101000110;
	 w_i = 24'b 111111111111111101010001;
	 next_valid = 1'b1;
	 end
	11'd1414: begin 
	 w_r = 24'b 111111111111111101000100;
	 w_i = 24'b 111111111111111101010010;
	 next_valid = 1'b1;
	 end
	11'd1415: begin 
	 w_r = 24'b 111111111111111101000011;
	 w_i = 24'b 111111111111111101010011;
	 next_valid = 1'b1;
	 end
	11'd1416: begin 
	 w_r = 24'b 111111111111111101000010;
	 w_i = 24'b 111111111111111101010100;
	 next_valid = 1'b1;
	 end
	11'd1417: begin 
	 w_r = 24'b 111111111111111101000001;
	 w_i = 24'b 111111111111111101010101;
	 next_valid = 1'b1;
	 end
	11'd1418: begin 
	 w_r = 24'b 111111111111111101000000;
	 w_i = 24'b 111111111111111101010110;
	 next_valid = 1'b1;
	 end
	11'd1419: begin 
	 w_r = 24'b 111111111111111100111111;
	 w_i = 24'b 111111111111111101011000;
	 next_valid = 1'b1;
	 end
	11'd1420: begin 
	 w_r = 24'b 111111111111111100111110;
	 w_i = 24'b 111111111111111101011001;
	 next_valid = 1'b1;
	 end
	11'd1421: begin 
	 w_r = 24'b 111111111111111100111101;
	 w_i = 24'b 111111111111111101011010;
	 next_valid = 1'b1;
	 end
	11'd1422: begin 
	 w_r = 24'b 111111111111111100111100;
	 w_i = 24'b 111111111111111101011011;
	 next_valid = 1'b1;
	 end
	11'd1423: begin 
	 w_r = 24'b 111111111111111100111011;
	 w_i = 24'b 111111111111111101011100;
	 next_valid = 1'b1;
	 end
	11'd1424: begin 
	 w_r = 24'b 111111111111111100111010;
	 w_i = 24'b 111111111111111101011110;
	 next_valid = 1'b1;
	 end
	11'd1425: begin 
	 w_r = 24'b 111111111111111100111001;
	 w_i = 24'b 111111111111111101011111;
	 next_valid = 1'b1;
	 end
	11'd1426: begin 
	 w_r = 24'b 111111111111111100111000;
	 w_i = 24'b 111111111111111101100000;
	 next_valid = 1'b1;
	 end
	11'd1427: begin 
	 w_r = 24'b 111111111111111100110111;
	 w_i = 24'b 111111111111111101100001;
	 next_valid = 1'b1;
	 end
	11'd1428: begin 
	 w_r = 24'b 111111111111111100110110;
	 w_i = 24'b 111111111111111101100011;
	 next_valid = 1'b1;
	 end
	11'd1429: begin 
	 w_r = 24'b 111111111111111100110101;
	 w_i = 24'b 111111111111111101100100;
	 next_valid = 1'b1;
	 end
	11'd1430: begin 
	 w_r = 24'b 111111111111111100110100;
	 w_i = 24'b 111111111111111101100101;
	 next_valid = 1'b1;
	 end
	11'd1431: begin 
	 w_r = 24'b 111111111111111100110011;
	 w_i = 24'b 111111111111111101100110;
	 next_valid = 1'b1;
	 end
	11'd1432: begin 
	 w_r = 24'b 111111111111111100110010;
	 w_i = 24'b 111111111111111101101000;
	 next_valid = 1'b1;
	 end
	11'd1433: begin 
	 w_r = 24'b 111111111111111100110001;
	 w_i = 24'b 111111111111111101101001;
	 next_valid = 1'b1;
	 end
	11'd1434: begin 
	 w_r = 24'b 111111111111111100110001;
	 w_i = 24'b 111111111111111101101010;
	 next_valid = 1'b1;
	 end
	11'd1435: begin 
	 w_r = 24'b 111111111111111100110000;
	 w_i = 24'b 111111111111111101101011;
	 next_valid = 1'b1;
	 end
	11'd1436: begin 
	 w_r = 24'b 111111111111111100101111;
	 w_i = 24'b 111111111111111101101101;
	 next_valid = 1'b1;
	 end
	11'd1437: begin 
	 w_r = 24'b 111111111111111100101110;
	 w_i = 24'b 111111111111111101101110;
	 next_valid = 1'b1;
	 end
	11'd1438: begin 
	 w_r = 24'b 111111111111111100101101;
	 w_i = 24'b 111111111111111101101111;
	 next_valid = 1'b1;
	 end
	11'd1439: begin 
	 w_r = 24'b 111111111111111100101100;
	 w_i = 24'b 111111111111111101110000;
	 next_valid = 1'b1;
	 end
	11'd1440: begin 
	 w_r = 24'b 111111111111111100101011;
	 w_i = 24'b 111111111111111101110010;
	 next_valid = 1'b1;
	 end
	11'd1441: begin 
	 w_r = 24'b 111111111111111100101010;
	 w_i = 24'b 111111111111111101110011;
	 next_valid = 1'b1;
	 end
	11'd1442: begin 
	 w_r = 24'b 111111111111111100101001;
	 w_i = 24'b 111111111111111101110100;
	 next_valid = 1'b1;
	 end
	11'd1443: begin 
	 w_r = 24'b 111111111111111100101001;
	 w_i = 24'b 111111111111111101110110;
	 next_valid = 1'b1;
	 end
	11'd1444: begin 
	 w_r = 24'b 111111111111111100101000;
	 w_i = 24'b 111111111111111101110111;
	 next_valid = 1'b1;
	 end
	11'd1445: begin 
	 w_r = 24'b 111111111111111100100111;
	 w_i = 24'b 111111111111111101111000;
	 next_valid = 1'b1;
	 end
	11'd1446: begin 
	 w_r = 24'b 111111111111111100100110;
	 w_i = 24'b 111111111111111101111010;
	 next_valid = 1'b1;
	 end
	11'd1447: begin 
	 w_r = 24'b 111111111111111100100101;
	 w_i = 24'b 111111111111111101111011;
	 next_valid = 1'b1;
	 end
	11'd1448: begin 
	 w_r = 24'b 111111111111111100100100;
	 w_i = 24'b 111111111111111101111100;
	 next_valid = 1'b1;
	 end
	11'd1449: begin 
	 w_r = 24'b 111111111111111100100100;
	 w_i = 24'b 111111111111111101111110;
	 next_valid = 1'b1;
	 end
	11'd1450: begin 
	 w_r = 24'b 111111111111111100100011;
	 w_i = 24'b 111111111111111101111111;
	 next_valid = 1'b1;
	 end
	11'd1451: begin 
	 w_r = 24'b 111111111111111100100010;
	 w_i = 24'b 111111111111111110000000;
	 next_valid = 1'b1;
	 end
	11'd1452: begin 
	 w_r = 24'b 111111111111111100100001;
	 w_i = 24'b 111111111111111110000010;
	 next_valid = 1'b1;
	 end
	11'd1453: begin 
	 w_r = 24'b 111111111111111100100000;
	 w_i = 24'b 111111111111111110000011;
	 next_valid = 1'b1;
	 end
	11'd1454: begin 
	 w_r = 24'b 111111111111111100100000;
	 w_i = 24'b 111111111111111110000101;
	 next_valid = 1'b1;
	 end
	11'd1455: begin 
	 w_r = 24'b 111111111111111100011111;
	 w_i = 24'b 111111111111111110000110;
	 next_valid = 1'b1;
	 end
	11'd1456: begin 
	 w_r = 24'b 111111111111111100011110;
	 w_i = 24'b 111111111111111110000111;
	 next_valid = 1'b1;
	 end
	11'd1457: begin 
	 w_r = 24'b 111111111111111100011101;
	 w_i = 24'b 111111111111111110001001;
	 next_valid = 1'b1;
	 end
	11'd1458: begin 
	 w_r = 24'b 111111111111111100011101;
	 w_i = 24'b 111111111111111110001010;
	 next_valid = 1'b1;
	 end
	11'd1459: begin 
	 w_r = 24'b 111111111111111100011100;
	 w_i = 24'b 111111111111111110001011;
	 next_valid = 1'b1;
	 end
	11'd1460: begin 
	 w_r = 24'b 111111111111111100011011;
	 w_i = 24'b 111111111111111110001101;
	 next_valid = 1'b1;
	 end
	11'd1461: begin 
	 w_r = 24'b 111111111111111100011011;
	 w_i = 24'b 111111111111111110001110;
	 next_valid = 1'b1;
	 end
	11'd1462: begin 
	 w_r = 24'b 111111111111111100011010;
	 w_i = 24'b 111111111111111110010000;
	 next_valid = 1'b1;
	 end
	11'd1463: begin 
	 w_r = 24'b 111111111111111100011001;
	 w_i = 24'b 111111111111111110010001;
	 next_valid = 1'b1;
	 end
	11'd1464: begin 
	 w_r = 24'b 111111111111111100011001;
	 w_i = 24'b 111111111111111110010011;
	 next_valid = 1'b1;
	 end
	11'd1465: begin 
	 w_r = 24'b 111111111111111100011000;
	 w_i = 24'b 111111111111111110010100;
	 next_valid = 1'b1;
	 end
	11'd1466: begin 
	 w_r = 24'b 111111111111111100010111;
	 w_i = 24'b 111111111111111110010101;
	 next_valid = 1'b1;
	 end
	11'd1467: begin 
	 w_r = 24'b 111111111111111100010111;
	 w_i = 24'b 111111111111111110010111;
	 next_valid = 1'b1;
	 end
	11'd1468: begin 
	 w_r = 24'b 111111111111111100010110;
	 w_i = 24'b 111111111111111110011000;
	 next_valid = 1'b1;
	 end
	11'd1469: begin 
	 w_r = 24'b 111111111111111100010101;
	 w_i = 24'b 111111111111111110011010;
	 next_valid = 1'b1;
	 end
	11'd1470: begin 
	 w_r = 24'b 111111111111111100010101;
	 w_i = 24'b 111111111111111110011011;
	 next_valid = 1'b1;
	 end
	11'd1471: begin 
	 w_r = 24'b 111111111111111100010100;
	 w_i = 24'b 111111111111111110011101;
	 next_valid = 1'b1;
	 end
	11'd1472: begin 
	 w_r = 24'b 111111111111111100010011;
	 w_i = 24'b 111111111111111110011110;
	 next_valid = 1'b1;
	 end
	11'd1473: begin 
	 w_r = 24'b 111111111111111100010011;
	 w_i = 24'b 111111111111111110011111;
	 next_valid = 1'b1;
	 end
	11'd1474: begin 
	 w_r = 24'b 111111111111111100010010;
	 w_i = 24'b 111111111111111110100001;
	 next_valid = 1'b1;
	 end
	11'd1475: begin 
	 w_r = 24'b 111111111111111100010010;
	 w_i = 24'b 111111111111111110100010;
	 next_valid = 1'b1;
	 end
	11'd1476: begin 
	 w_r = 24'b 111111111111111100010001;
	 w_i = 24'b 111111111111111110100100;
	 next_valid = 1'b1;
	 end
	11'd1477: begin 
	 w_r = 24'b 111111111111111100010001;
	 w_i = 24'b 111111111111111110100101;
	 next_valid = 1'b1;
	 end
	11'd1478: begin 
	 w_r = 24'b 111111111111111100010000;
	 w_i = 24'b 111111111111111110100111;
	 next_valid = 1'b1;
	 end
	11'd1479: begin 
	 w_r = 24'b 111111111111111100001111;
	 w_i = 24'b 111111111111111110101000;
	 next_valid = 1'b1;
	 end
	11'd1480: begin 
	 w_r = 24'b 111111111111111100001111;
	 w_i = 24'b 111111111111111110101010;
	 next_valid = 1'b1;
	 end
	11'd1481: begin 
	 w_r = 24'b 111111111111111100001110;
	 w_i = 24'b 111111111111111110101011;
	 next_valid = 1'b1;
	 end
	11'd1482: begin 
	 w_r = 24'b 111111111111111100001110;
	 w_i = 24'b 111111111111111110101101;
	 next_valid = 1'b1;
	 end
	11'd1483: begin 
	 w_r = 24'b 111111111111111100001101;
	 w_i = 24'b 111111111111111110101110;
	 next_valid = 1'b1;
	 end
	11'd1484: begin 
	 w_r = 24'b 111111111111111100001101;
	 w_i = 24'b 111111111111111110110000;
	 next_valid = 1'b1;
	 end
	11'd1485: begin 
	 w_r = 24'b 111111111111111100001100;
	 w_i = 24'b 111111111111111110110001;
	 next_valid = 1'b1;
	 end
	11'd1486: begin 
	 w_r = 24'b 111111111111111100001100;
	 w_i = 24'b 111111111111111110110011;
	 next_valid = 1'b1;
	 end
	11'd1487: begin 
	 w_r = 24'b 111111111111111100001011;
	 w_i = 24'b 111111111111111110110100;
	 next_valid = 1'b1;
	 end
	11'd1488: begin 
	 w_r = 24'b 111111111111111100001011;
	 w_i = 24'b 111111111111111110110110;
	 next_valid = 1'b1;
	 end
	11'd1489: begin 
	 w_r = 24'b 111111111111111100001011;
	 w_i = 24'b 111111111111111110110111;
	 next_valid = 1'b1;
	 end
	11'd1490: begin 
	 w_r = 24'b 111111111111111100001010;
	 w_i = 24'b 111111111111111110111001;
	 next_valid = 1'b1;
	 end
	11'd1491: begin 
	 w_r = 24'b 111111111111111100001010;
	 w_i = 24'b 111111111111111110111010;
	 next_valid = 1'b1;
	 end
	11'd1492: begin 
	 w_r = 24'b 111111111111111100001001;
	 w_i = 24'b 111111111111111110111100;
	 next_valid = 1'b1;
	 end
	11'd1493: begin 
	 w_r = 24'b 111111111111111100001001;
	 w_i = 24'b 111111111111111110111101;
	 next_valid = 1'b1;
	 end
	11'd1494: begin 
	 w_r = 24'b 111111111111111100001000;
	 w_i = 24'b 111111111111111110111111;
	 next_valid = 1'b1;
	 end
	11'd1495: begin 
	 w_r = 24'b 111111111111111100001000;
	 w_i = 24'b 111111111111111111000000;
	 next_valid = 1'b1;
	 end
	11'd1496: begin 
	 w_r = 24'b 111111111111111100001000;
	 w_i = 24'b 111111111111111111000010;
	 next_valid = 1'b1;
	 end
	11'd1497: begin 
	 w_r = 24'b 111111111111111100000111;
	 w_i = 24'b 111111111111111111000011;
	 next_valid = 1'b1;
	 end
	11'd1498: begin 
	 w_r = 24'b 111111111111111100000111;
	 w_i = 24'b 111111111111111111000101;
	 next_valid = 1'b1;
	 end
	11'd1499: begin 
	 w_r = 24'b 111111111111111100000111;
	 w_i = 24'b 111111111111111111000110;
	 next_valid = 1'b1;
	 end
	11'd1500: begin 
	 w_r = 24'b 111111111111111100000110;
	 w_i = 24'b 111111111111111111001000;
	 next_valid = 1'b1;
	 end
	11'd1501: begin 
	 w_r = 24'b 111111111111111100000110;
	 w_i = 24'b 111111111111111111001001;
	 next_valid = 1'b1;
	 end
	11'd1502: begin 
	 w_r = 24'b 111111111111111100000110;
	 w_i = 24'b 111111111111111111001011;
	 next_valid = 1'b1;
	 end
	11'd1503: begin 
	 w_r = 24'b 111111111111111100000101;
	 w_i = 24'b 111111111111111111001101;
	 next_valid = 1'b1;
	 end
	11'd1504: begin 
	 w_r = 24'b 111111111111111100000101;
	 w_i = 24'b 111111111111111111001110;
	 next_valid = 1'b1;
	 end
	11'd1505: begin 
	 w_r = 24'b 111111111111111100000101;
	 w_i = 24'b 111111111111111111010000;
	 next_valid = 1'b1;
	 end
	11'd1506: begin 
	 w_r = 24'b 111111111111111100000100;
	 w_i = 24'b 111111111111111111010001;
	 next_valid = 1'b1;
	 end
	11'd1507: begin 
	 w_r = 24'b 111111111111111100000100;
	 w_i = 24'b 111111111111111111010011;
	 next_valid = 1'b1;
	 end
	11'd1508: begin 
	 w_r = 24'b 111111111111111100000100;
	 w_i = 24'b 111111111111111111010100;
	 next_valid = 1'b1;
	 end
	11'd1509: begin 
	 w_r = 24'b 111111111111111100000100;
	 w_i = 24'b 111111111111111111010110;
	 next_valid = 1'b1;
	 end
	11'd1510: begin 
	 w_r = 24'b 111111111111111100000011;
	 w_i = 24'b 111111111111111111010111;
	 next_valid = 1'b1;
	 end
	11'd1511: begin 
	 w_r = 24'b 111111111111111100000011;
	 w_i = 24'b 111111111111111111011001;
	 next_valid = 1'b1;
	 end
	11'd1512: begin 
	 w_r = 24'b 111111111111111100000011;
	 w_i = 24'b 111111111111111111011010;
	 next_valid = 1'b1;
	 end
	11'd1513: begin 
	 w_r = 24'b 111111111111111100000011;
	 w_i = 24'b 111111111111111111011100;
	 next_valid = 1'b1;
	 end
	11'd1514: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111011110;
	 next_valid = 1'b1;
	 end
	11'd1515: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111011111;
	 next_valid = 1'b1;
	 end
	11'd1516: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111100001;
	 next_valid = 1'b1;
	 end
	11'd1517: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111100010;
	 next_valid = 1'b1;
	 end
	11'd1518: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111100100;
	 next_valid = 1'b1;
	 end
	11'd1519: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111100101;
	 next_valid = 1'b1;
	 end
	11'd1520: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111100111;
	 next_valid = 1'b1;
	 end
	11'd1521: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111101000;
	 next_valid = 1'b1;
	 end
	11'd1522: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111101010;
	 next_valid = 1'b1;
	 end
	11'd1523: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111101100;
	 next_valid = 1'b1;
	 end
	11'd1524: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111101101;
	 next_valid = 1'b1;
	 end
	11'd1525: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111101111;
	 next_valid = 1'b1;
	 end
	11'd1526: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110000;
	 next_valid = 1'b1;
	 end
	11'd1527: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110010;
	 next_valid = 1'b1;
	 end
	11'd1528: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110011;
	 next_valid = 1'b1;
	 end
	11'd1529: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110101;
	 next_valid = 1'b1;
	 end
	11'd1530: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110111;
	 next_valid = 1'b1;
	 end
	11'd1531: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111111000;
	 next_valid = 1'b1;
	 end
	11'd1532: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111111010;
	 next_valid = 1'b1;
	 end
	11'd1533: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111111011;
	 next_valid = 1'b1;
	 end
	11'd1534: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111111101;
	 next_valid = 1'b1;
	 end
	11'd1535: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111111110;
	 next_valid = 1'b0;
	 end
	default: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 000000000000000000000000;
	 next_valid = 1'b1;
	 end
	endcase

end

always@(posedge clk or negedge rst_n)begin
    if(~rst_n)begin
        count <= 0;
        valid <= 0;
    end
    else if(in_valid)
    begin
        count <= next_count;
        valid <= in_valid;
    end
    else if (valid)
    begin
        count <= next_count;
        valid <= next_valid;
    end
end
endmodule