module FFT(
input clk,
input rst_n,
input in_valid,
input signed [11:0] din_r,
input signed [11:0] din_i,
output out_valid,
output reg signed [15:0] dout_r,
output reg signed [15:0] dout_i
);
//////////////////////////////////////////////////////////////
// Declaration:
integer i;
reg signed  [15:0] result_r[0:1023];
reg signed  [15:0] result_i[0:1023];
reg signed  [15:0] result_r_ns[0:1023];
reg signed  [15:0] result_i_ns[0:1023];
reg signed [15:0] next_dout_r;
reg signed [15:0] next_dout_i;
reg         [10:0]   count_y;
reg         [10:0]   next_count_y;

reg signed [23:0] din_r_reg,din_i_reg;
reg in_valid_reg,r9_valid,next_r9_valid;
reg [1:0] no10_state;
reg s10_count,next_s10_count;
reg next_over,over;
reg assign_out;
reg next_out_valid;
reg [9:0]y_1_delay;

wire [23:0] out_r,out_i;
wire [9:0] y_1;
wire [23:0] din_r_wire,din_i_wire;

assign out_valid = assign_out;
assign y_1 = (count_y>10'd0)? (count_y - 10'd1) : count_y; 
assign din_r_wire = din_r_reg;
assign din_i_wire = din_i_reg;

wire [1:0] rom512_state;
wire [23:0]rom512_w_r,rom512_w_i;
wire [23:0]shift_512_dout_r,shift_512_dout_i;
wire [23:0]radix_no1_op_r,radix_no1_op_i;
wire [23:0]radix_no1_delay_r,radix_no1_delay_i;
wire radix_no1_outvalid;

wire [1:0] rom256_state;
wire [23:0]rom256_w_r,rom256_w_i;
wire [23:0]shift_256_dout_r,shift_256_dout_i;
wire [23:0]radix_no2_delay_r,radix_no2_delay_i;
wire [23:0]radix_no2_op_r,radix_no2_op_i;
wire radix_no2_outvalid;

wire [1:0] rom128_state;
wire [23:0]rom128_w_r,rom128_w_i;
wire [23:0]shift_128_dout_r,shift_128_dout_i;
wire [23:0]radix_no3_delay_r,radix_no3_delay_i;
wire [23:0]radix_no3_op_r,radix_no3_op_i;
wire radix_no3_outvalid;

wire [1:0] rom64_state;
wire [23:0]rom64_w_r,rom64_w_i;
wire [23:0]shift_64_dout_r,shift_64_dout_i;
wire [23:0]radix_no4_delay_r,radix_no4_delay_i;
wire [23:0]radix_no4_op_r,radix_no4_op_i;
wire radix_no4_outvalid;

wire [1:0] rom32_state;
wire [23:0]rom32_w_r,rom32_w_i;
wire [23:0]shift_32_dout_r,shift_32_dout_i;
wire [23:0]radix_no5_delay_r,radix_no5_delay_i;
wire [23:0]radix_no5_op_r,radix_no5_op_i;
wire radix_no5_outvalid;

wire [1:0] rom16_state;
wire [23:0]rom16_w_r,rom16_w_i;
wire [23:0]shift_16_dout_r,shift_16_dout_i;
wire [23:0]radix_no6_delay_r,radix_no6_delay_i;
wire [23:0]radix_no6_op_r,radix_no6_op_i;
wire radix_no6_outvalid;

wire [1:0] rom8_state;
wire [23:0]rom8_w_r,rom8_w_i;
wire [23:0]shift_8_dout_r,shift_8_dout_i;
wire [23:0]radix_no7_delay_r,radix_no7_delay_i;
wire [23:0]radix_no7_op_r,radix_no7_op_i;
wire radix_no7_outvalid;

wire [1:0] rom4_state;
wire [23:0]rom4_w_r,rom4_w_i;
wire [23:0]shift_4_dout_r,shift_4_dout_i;
wire [23:0]radix_no8_delay_r,radix_no8_delay_i;
wire [23:0]radix_no8_op_r,radix_no8_op_i;
wire radix_no8_outvalid;

wire [1:0] rom2_state;
wire [23:0]rom2_w_r,rom2_w_i;
wire [23:0]shift_2_dout_r,shift_2_dout_i;
wire [23:0]radix_no9_delay_r,radix_no9_delay_i;
wire [23:0]radix_no9_op_r,radix_no9_op_i;
wire radix_no9_outvalid;

wire [23:0]shift_1_dout_r,shift_1_dout_i;
wire [23:0]radix_no10_delay_r,radix_no10_delay_i;
wire [23:0]radix_no10_op_r,radix_no10_op_i;

//////////////////////////////////////////////////////////////
// Step 1:
radix2 radix_no1(
.state(rom512_state),//state ctrl
.din_a_r(shift_512_dout_r),//fb
.din_a_i(shift_512_dout_i),//fb
.din_b_r(din_r_wire),//input
.din_b_i(din_i_wire),//input
.w_r(rom512_w_r),//twindle_r
.w_i(rom512_w_i),//twindle_i
.op_r(radix_no1_op_r),
.op_i(radix_no1_op_i),
.delay_r(radix_no1_delay_r),
.delay_i(radix_no1_delay_i),
.outvalid(radix_no1_outvalid)
);

shift_512 shift_512(
.clk(clk),.rst_n(rst_n),
.in_valid(in_valid_reg),
.din_r(radix_no1_delay_r),
.din_i(radix_no1_delay_i),
.dout_r(shift_512_dout_r),
.dout_i(shift_512_dout_i)
);

ROM_512 rom512(
.clk(clk),
.in_valid(in_valid_reg),
.rst_n(rst_n),
.w_r(rom512_w_r),
.w_i(rom512_w_i),
.state(rom512_state)
);

// Step 2:
radix2 radix_no2(
.state(rom256_state),//state ctrl
.din_a_r(shift_256_dout_r),//fb
.din_a_i(shift_256_dout_i),//fb
.din_b_r(radix_no1_op_r),//input
.din_b_i(radix_no1_op_i),//input
.w_r(rom256_w_r),//twindle
.w_i(rom256_w_i),//d
.op_r(radix_no2_op_r),
.op_i(radix_no2_op_i),
.delay_r(radix_no2_delay_r),
.delay_i(radix_no2_delay_i),
.outvalid(radix_no2_outvalid)
);

shift_256 shift_256(
.clk(clk),.rst_n(rst_n),
.in_valid(radix_no1_outvalid),
.din_r(radix_no2_delay_r),
.din_i(radix_no2_delay_i),
.dout_r(shift_256_dout_r),
.dout_i(shift_256_dout_i)
);

ROM_256 rom256(
.clk(clk),
.in_valid(radix_no1_outvalid),
.rst_n(rst_n),
.w_r(rom256_w_r),
.w_i(rom256_w_i),
.state(rom256_state)
);

// Step 3:
radix2 radix_no3(
.state(rom128_state),//state ctrl
.din_a_r(shift_128_dout_r),//fb
.din_a_i(shift_128_dout_i),//fb
.din_b_r(radix_no2_op_r),//input
.din_b_i(radix_no2_op_i),//input
.w_r(rom128_w_r),//twindle
.w_i(rom128_w_i),//d
.op_r(radix_no3_op_r),
.op_i(radix_no3_op_i),
.delay_r(radix_no3_delay_r),
.delay_i(radix_no3_delay_i),
.outvalid(radix_no3_outvalid)
);

shift_128 shift_128(
.clk(clk),.rst_n(rst_n),
.in_valid(radix_no2_outvalid),
.din_r(radix_no3_delay_r),
.din_i(radix_no3_delay_i),
.dout_r(shift_128_dout_r),
.dout_i(shift_128_dout_i)  
);

ROM_128 rom128(
.clk(clk),
.in_valid(radix_no2_outvalid),
.rst_n(rst_n),
.w_r(rom128_w_r),
.w_i(rom128_w_i),
.state(rom128_state)
);

// Step 4:
radix2 radix_no4(
.state(rom64_state),//state ctrl
.din_a_r(shift_64_dout_r),//fb
.din_a_i(shift_64_dout_i),//fb
.din_b_r(radix_no3_op_r),//input
.din_b_i(radix_no3_op_i),//input
.w_r(rom64_w_r),//twindle
.w_i(rom64_w_i),//d
.op_r(radix_no4_op_r),
.op_i(radix_no4_op_i),
.delay_r(radix_no4_delay_r),
.delay_i(radix_no4_delay_i),
.outvalid(radix_no4_outvalid)
);

shift_64 shift_64(
.clk(clk),.rst_n(rst_n),
.in_valid(radix_no3_outvalid),
.din_r(radix_no4_delay_r),
.din_i(radix_no4_delay_i),
.dout_r(shift_64_dout_r),
.dout_i(shift_64_dout_i)
);

ROM_64 rom64(
.clk(clk),
.in_valid(radix_no3_outvalid),
.rst_n(rst_n),
.w_r(rom64_w_r),
.w_i(rom64_w_i),
.state(rom64_state)
);

// Step 5:
radix2 radix_no5(
.state(rom32_state),//state ctrl
.din_a_r(shift_32_dout_r),//fb
.din_a_i(shift_32_dout_i),//fb
.din_b_r(radix_no4_op_r),//input
.din_b_i(radix_no4_op_i),//input
.w_r(rom32_w_r),//twindle
.w_i(rom32_w_i),//d
.op_r(radix_no5_op_r),
.op_i(radix_no5_op_i),
.delay_r(radix_no5_delay_r),
.delay_i(radix_no5_delay_i),
.outvalid(radix_no5_outvalid)
);

shift_32 shift_32(
.clk(clk),.rst_n(rst_n),
.in_valid(radix_no4_outvalid),
.din_r(radix_no5_delay_r),
.din_i(radix_no5_delay_i),
.dout_r(shift_32_dout_r),
.dout_i(shift_32_dout_i)
);

ROM_32 rom32(
.clk(clk),
.in_valid(radix_no4_outvalid),
.rst_n(rst_n),
.w_r(rom32_w_r),
.w_i(rom32_w_i),
.state(rom32_state)
);

// Step 6:
radix2 radix_no6(
.state(rom16_state),//state ctrl
.din_a_r(shift_16_dout_r),//fb
.din_a_i(shift_16_dout_i),//fb
.din_b_r(radix_no5_op_r),//input
.din_b_i(radix_no5_op_i),//input
.w_r(rom16_w_r),//twindle
.w_i(rom16_w_i),//d
.op_r(radix_no6_op_r),
.op_i(radix_no6_op_i),
.delay_r(radix_no6_delay_r),
.delay_i(radix_no6_delay_i),
.outvalid(radix_no6_outvalid)
);

shift_16 shift_16(
.clk(clk),.rst_n(rst_n),
.in_valid(radix_no5_outvalid),
.din_r(radix_no6_delay_r),
.din_i(radix_no6_delay_i),
.dout_r(shift_16_dout_r),
.dout_i(shift_16_dout_i)
);

ROM_16 rom16(
.clk(clk),
.in_valid(radix_no5_outvalid),
.rst_n(rst_n),
.w_r(rom16_w_r),
.w_i(rom16_w_i),
.state(rom16_state)
);

// Step 7:
radix2 radix_no7(
.state(rom8_state),//state ctrl
.din_a_r(shift_8_dout_r),//fb
.din_a_i(shift_8_dout_i),//fb
.din_b_r(radix_no6_op_r),//input
.din_b_i(radix_no6_op_i),//input
.w_r(rom8_w_r),//twindle
.w_i(rom8_w_i),//d
.op_r(radix_no7_op_r),
.op_i(radix_no7_op_i),
.delay_r(radix_no7_delay_r),
.delay_i(radix_no7_delay_i),
.outvalid(radix_no7_outvalid)
);

shift_8 shift_8(
.clk(clk),.rst_n(rst_n),
.in_valid(radix_no6_outvalid),
.din_r(radix_no7_delay_r),
.din_i(radix_no7_delay_i),
.dout_r(shift_8_dout_r),
.dout_i(shift_8_dout_i)
);

ROM_8 rom8(
.clk(clk),
.in_valid(radix_no6_outvalid),
.rst_n(rst_n),
.w_r(rom8_w_r),
.w_i(rom8_w_i),
.state(rom8_state)
);

// Step 8:
radix2 radix_no8(
.state(rom4_state),//state ctrl
.din_a_r(shift_4_dout_r),//fb
.din_a_i(shift_4_dout_i),//fb
.din_b_r(radix_no7_op_r),//input
.din_b_i(radix_no7_op_i),//input
.w_r(rom4_w_r),//twindle
.w_i(rom4_w_i),//d
.op_r(radix_no8_op_r),
.op_i(radix_no8_op_i),
.delay_r(radix_no8_delay_r),
.delay_i(radix_no8_delay_i),
.outvalid(radix_no8_outvalid)
);

shift_4 shift_4(
.clk(clk),.rst_n(rst_n),
.in_valid(radix_no7_outvalid),
.din_r(radix_no8_delay_r),
.din_i(radix_no8_delay_i),
.dout_r(shift_4_dout_r),
.dout_i(shift_4_dout_i)
);

ROM_4 rom4(
.clk(clk),
.in_valid(radix_no7_outvalid),
.rst_n(rst_n),
.w_r(rom4_w_r),
.w_i(rom4_w_i),
.state(rom4_state)
);

// Step 9:
radix2 radix_no9(
.state(rom2_state),//state ctrl
.din_a_r(shift_2_dout_r),//fb
.din_a_i(shift_2_dout_i),//fb
.din_b_r(radix_no8_op_r),//input
.din_b_i(radix_no8_op_i),//input
.w_r(rom2_w_r),//twindle
.w_i(rom2_w_i),//d
.op_r(radix_no9_op_r),
.op_i(radix_no9_op_i),
.delay_r(radix_no9_delay_r),
.delay_i(radix_no9_delay_i),
.outvalid(radix_no9_outvalid)
);

shift_2 shift_2(
.clk(clk),.rst_n(rst_n),
.in_valid(radix_no8_outvalid),
.din_r(radix_no9_delay_r),
.din_i(radix_no9_delay_i),
.dout_r(shift_2_dout_r),
.dout_i(shift_2_dout_i)
);

ROM_2 rom2(
.clk(clk),
.in_valid(radix_no8_outvalid),
.rst_n(rst_n),
.w_r(rom2_w_r),
.w_i(rom2_w_i),
.state(rom2_state)
);

// Step 10:
radix2 radix_no10(
.state(no10_state),//state ctrl
.din_a_r(shift_1_dout_r),//fb
.din_a_i(shift_1_dout_i),//fb
.din_b_r(radix_no9_op_r),//input
.din_b_i(radix_no9_op_i),//input
.w_r(24'd256),//twindle
.w_i(24'd0),//d
.op_r(out_r),
.op_i(out_i),
.delay_r(radix_no10_delay_r),
.delay_i(radix_no10_delay_i),
.outvalid()
);

shift_1 shift_1(
.clk(clk),.rst_n(rst_n),
.in_valid(radix_no9_outvalid),
.din_r(radix_no10_delay_r),
.din_i(radix_no10_delay_i),
.dout_r(shift_1_dout_r),
.dout_i(shift_1_dout_i)
);

//////////////////////////////////////////////////////////////
always@(*)begin

    next_r9_valid = radix_no9_outvalid;
    if (r9_valid)next_s10_count = s10_count + 1;
    else next_s10_count = s10_count;
    
    if(r9_valid && s10_count == 1'b0)no10_state = 2'b01;
    else if(r9_valid && s10_count == 1'b1)no10_state = 2'b10;
    else no10_state = 2'b00;

    if(radix_no9_outvalid) next_count_y = count_y + 10'd1;
    else next_count_y = count_y;

    if(next_out_valid) begin
        next_dout_r = result_r[y_1_delay];
        next_dout_i = result_i[y_1_delay];
    end
    else begin
        next_dout_r = dout_r;
        next_dout_i = dout_i;
    end
end
//////////////////////////////////////////////////////////////
always@(posedge clk or negedge rst_n)begin
    if(~rst_n)begin
        din_r_reg <= 0;
        din_i_reg <= 0;
        in_valid_reg <= 0;
        s10_count <= 0;
        r9_valid <= 0;
        count_y <= 0;
        assign_out <= 0;
        over <= 0;
        dout_r <= 0;
        dout_i <= 0;
        y_1_delay <= 0;
        for (i=0;i<=1023;i=i+1) begin
            result_r[i] <= 0;
            result_i[i] <= 0;
        end
    end
    else begin
        din_r_reg <= {{4{din_r[11]}},din_r,8'b0};
        din_i_reg <= {{4{din_i[11]}},din_i,8'b0};
        in_valid_reg <= in_valid;
        s10_count <= next_s10_count;
        r9_valid <= next_r9_valid;
        count_y  <= next_count_y;
        assign_out <= next_out_valid;
        over <= next_over;
        y_1_delay <= y_1;
        dout_r <= next_dout_r;
        dout_i <= next_dout_i;
        for (i=0;i<=1023;i=i+1) begin
            result_r[i] <= result_r_ns[i];
            result_i[i] <= result_i_ns[i];
        end
    end
end
//////////////////////////////////////////////////////////////
// Sorting module:
always @(*) begin

    next_over = over;
    for (i=0;i<=1023;i=i+1) begin
        result_r_ns[i] = result_r[i];
        result_i_ns[i] = result_i[i];
    end
    if(next_over==1'b1)next_out_valid = 1'b1;
    else next_out_valid = assign_out;

    if(over!=1'b1) begin
        case((y_1))
        10'd0 : begin
           result_r_ns[1023] = out_r[23:8];
           result_i_ns[1023] = out_i[23:8];
        end
        10'd1 : begin
           result_r_ns[511] = out_r[23:8];
           result_i_ns[511] = out_i[23:8];
        end
        10'd2 : begin
           result_r_ns[255] = out_r[23:8];
           result_i_ns[255] = out_i[23:8];
        end
        10'd3 : begin
           result_r_ns[767] = out_r[23:8];
           result_i_ns[767] = out_i[23:8];
        end
        10'd4 : begin
           result_r_ns[127] = out_r[23:8];
           result_i_ns[127] = out_i[23:8];
        end
        10'd5 : begin
           result_r_ns[639] = out_r[23:8];
           result_i_ns[639] = out_i[23:8];
        end
        10'd6 : begin
           result_r_ns[383] = out_r[23:8];
           result_i_ns[383] = out_i[23:8];
        end
        10'd7 : begin
           result_r_ns[895] = out_r[23:8];
           result_i_ns[895] = out_i[23:8];
        end
        10'd8 : begin
           result_r_ns[63] = out_r[23:8];
           result_i_ns[63] = out_i[23:8];
        end
        10'd9 : begin
           result_r_ns[575] = out_r[23:8];
           result_i_ns[575] = out_i[23:8];
        end
        10'd10 : begin
           result_r_ns[319] = out_r[23:8];
           result_i_ns[319] = out_i[23:8];
        end
        10'd11 : begin
           result_r_ns[831] = out_r[23:8];
           result_i_ns[831] = out_i[23:8];
        end
        10'd12 : begin
           result_r_ns[191] = out_r[23:8];
           result_i_ns[191] = out_i[23:8];
        end
        10'd13 : begin
           result_r_ns[703] = out_r[23:8];
           result_i_ns[703] = out_i[23:8];
        end
        10'd14 : begin
           result_r_ns[447] = out_r[23:8];
           result_i_ns[447] = out_i[23:8];
        end
        10'd15 : begin
           result_r_ns[959] = out_r[23:8];
           result_i_ns[959] = out_i[23:8];
        end
        10'd16 : begin
           result_r_ns[31] = out_r[23:8];
           result_i_ns[31] = out_i[23:8];
        end
        10'd17 : begin
           result_r_ns[543] = out_r[23:8];
           result_i_ns[543] = out_i[23:8];
        end
        10'd18 : begin
           result_r_ns[287] = out_r[23:8];
           result_i_ns[287] = out_i[23:8];
        end
        10'd19 : begin
           result_r_ns[799] = out_r[23:8];
           result_i_ns[799] = out_i[23:8];
        end
        10'd20 : begin
           result_r_ns[159] = out_r[23:8];
           result_i_ns[159] = out_i[23:8];
        end
        10'd21 : begin
           result_r_ns[671] = out_r[23:8];
           result_i_ns[671] = out_i[23:8];
        end
        10'd22 : begin
           result_r_ns[415] = out_r[23:8];
           result_i_ns[415] = out_i[23:8];
        end
        10'd23 : begin
           result_r_ns[927] = out_r[23:8];
           result_i_ns[927] = out_i[23:8];
        end
        10'd24 : begin
           result_r_ns[95] = out_r[23:8];
           result_i_ns[95] = out_i[23:8];
        end
        10'd25 : begin
           result_r_ns[607] = out_r[23:8];
           result_i_ns[607] = out_i[23:8];
        end
        10'd26 : begin
           result_r_ns[351] = out_r[23:8];
           result_i_ns[351] = out_i[23:8];
        end
        10'd27 : begin
           result_r_ns[863] = out_r[23:8];
           result_i_ns[863] = out_i[23:8];
        end
        10'd28 : begin
           result_r_ns[223] = out_r[23:8];
           result_i_ns[223] = out_i[23:8];
        end
        10'd29 : begin
           result_r_ns[735] = out_r[23:8];
           result_i_ns[735] = out_i[23:8];
        end
        10'd30 : begin
           result_r_ns[479] = out_r[23:8];
           result_i_ns[479] = out_i[23:8];
        end
        10'd31 : begin
           result_r_ns[991] = out_r[23:8];
           result_i_ns[991] = out_i[23:8];
        end
        10'd32 : begin
           result_r_ns[15] = out_r[23:8];
           result_i_ns[15] = out_i[23:8];
        end
        10'd33 : begin
           result_r_ns[527] = out_r[23:8];
           result_i_ns[527] = out_i[23:8];
        end
        10'd34 : begin
           result_r_ns[271] = out_r[23:8];
           result_i_ns[271] = out_i[23:8];
        end
        10'd35 : begin
           result_r_ns[783] = out_r[23:8];
           result_i_ns[783] = out_i[23:8];
        end
        10'd36 : begin
           result_r_ns[143] = out_r[23:8];
           result_i_ns[143] = out_i[23:8];
        end
        10'd37 : begin
           result_r_ns[655] = out_r[23:8];
           result_i_ns[655] = out_i[23:8];
        end
        10'd38 : begin
           result_r_ns[399] = out_r[23:8];
           result_i_ns[399] = out_i[23:8];
        end
        10'd39 : begin
           result_r_ns[911] = out_r[23:8];
           result_i_ns[911] = out_i[23:8];
        end
        10'd40 : begin
           result_r_ns[79] = out_r[23:8];
           result_i_ns[79] = out_i[23:8];
        end
        10'd41 : begin
           result_r_ns[591] = out_r[23:8];
           result_i_ns[591] = out_i[23:8];
        end
        10'd42 : begin
           result_r_ns[335] = out_r[23:8];
           result_i_ns[335] = out_i[23:8];
        end
        10'd43 : begin
           result_r_ns[847] = out_r[23:8];
           result_i_ns[847] = out_i[23:8];
        end
        10'd44 : begin
           result_r_ns[207] = out_r[23:8];
           result_i_ns[207] = out_i[23:8];
        end
        10'd45 : begin
           result_r_ns[719] = out_r[23:8];
           result_i_ns[719] = out_i[23:8];
        end
        10'd46 : begin
           result_r_ns[463] = out_r[23:8];
           result_i_ns[463] = out_i[23:8];
        end
        10'd47 : begin
           result_r_ns[975] = out_r[23:8];
           result_i_ns[975] = out_i[23:8];
        end
        10'd48 : begin
           result_r_ns[47] = out_r[23:8];
           result_i_ns[47] = out_i[23:8];
        end
        10'd49 : begin
           result_r_ns[559] = out_r[23:8];
           result_i_ns[559] = out_i[23:8];
        end
        10'd50 : begin
           result_r_ns[303] = out_r[23:8];
           result_i_ns[303] = out_i[23:8];
        end
        10'd51 : begin
           result_r_ns[815] = out_r[23:8];
           result_i_ns[815] = out_i[23:8];
        end
        10'd52 : begin
           result_r_ns[175] = out_r[23:8];
           result_i_ns[175] = out_i[23:8];
        end
        10'd53 : begin
           result_r_ns[687] = out_r[23:8];
           result_i_ns[687] = out_i[23:8];
        end
        10'd54 : begin
           result_r_ns[431] = out_r[23:8];
           result_i_ns[431] = out_i[23:8];
        end
        10'd55 : begin
           result_r_ns[943] = out_r[23:8];
           result_i_ns[943] = out_i[23:8];
        end
        10'd56 : begin
           result_r_ns[111] = out_r[23:8];
           result_i_ns[111] = out_i[23:8];
        end
        10'd57 : begin
           result_r_ns[623] = out_r[23:8];
           result_i_ns[623] = out_i[23:8];
        end
        10'd58 : begin
           result_r_ns[367] = out_r[23:8];
           result_i_ns[367] = out_i[23:8];
        end
        10'd59 : begin
           result_r_ns[879] = out_r[23:8];
           result_i_ns[879] = out_i[23:8];
        end
        10'd60 : begin
           result_r_ns[239] = out_r[23:8];
           result_i_ns[239] = out_i[23:8];
        end
        10'd61 : begin
           result_r_ns[751] = out_r[23:8];
           result_i_ns[751] = out_i[23:8];
        end
        10'd62 : begin
           result_r_ns[495] = out_r[23:8];
           result_i_ns[495] = out_i[23:8];
        end
        10'd63 : begin
           result_r_ns[1007] = out_r[23:8];
           result_i_ns[1007] = out_i[23:8];
        end
        10'd64 : begin
           result_r_ns[7] = out_r[23:8];
           result_i_ns[7] = out_i[23:8];
        end
        10'd65 : begin
           result_r_ns[519] = out_r[23:8];
           result_i_ns[519] = out_i[23:8];
        end
        10'd66 : begin
           result_r_ns[263] = out_r[23:8];
           result_i_ns[263] = out_i[23:8];
        end
        10'd67 : begin
           result_r_ns[775] = out_r[23:8];
           result_i_ns[775] = out_i[23:8];
        end
        10'd68 : begin
           result_r_ns[135] = out_r[23:8];
           result_i_ns[135] = out_i[23:8];
        end
        10'd69 : begin
           result_r_ns[647] = out_r[23:8];
           result_i_ns[647] = out_i[23:8];
        end
        10'd70 : begin
           result_r_ns[391] = out_r[23:8];
           result_i_ns[391] = out_i[23:8];
        end
        10'd71 : begin
           result_r_ns[903] = out_r[23:8];
           result_i_ns[903] = out_i[23:8];
        end
        10'd72 : begin
           result_r_ns[71] = out_r[23:8];
           result_i_ns[71] = out_i[23:8];
        end
        10'd73 : begin
           result_r_ns[583] = out_r[23:8];
           result_i_ns[583] = out_i[23:8];
        end
        10'd74 : begin
           result_r_ns[327] = out_r[23:8];
           result_i_ns[327] = out_i[23:8];
        end
        10'd75 : begin
           result_r_ns[839] = out_r[23:8];
           result_i_ns[839] = out_i[23:8];
        end
        10'd76 : begin
           result_r_ns[199] = out_r[23:8];
           result_i_ns[199] = out_i[23:8];
        end
        10'd77 : begin
           result_r_ns[711] = out_r[23:8];
           result_i_ns[711] = out_i[23:8];
        end
        10'd78 : begin
           result_r_ns[455] = out_r[23:8];
           result_i_ns[455] = out_i[23:8];
        end
        10'd79 : begin
           result_r_ns[967] = out_r[23:8];
           result_i_ns[967] = out_i[23:8];
        end
        10'd80 : begin
           result_r_ns[39] = out_r[23:8];
           result_i_ns[39] = out_i[23:8];
        end
        10'd81 : begin
           result_r_ns[551] = out_r[23:8];
           result_i_ns[551] = out_i[23:8];
        end
        10'd82 : begin
           result_r_ns[295] = out_r[23:8];
           result_i_ns[295] = out_i[23:8];
        end
        10'd83 : begin
           result_r_ns[807] = out_r[23:8];
           result_i_ns[807] = out_i[23:8];
        end
        10'd84 : begin
           result_r_ns[167] = out_r[23:8];
           result_i_ns[167] = out_i[23:8];
        end
        10'd85 : begin
           result_r_ns[679] = out_r[23:8];
           result_i_ns[679] = out_i[23:8];
        end
        10'd86 : begin
           result_r_ns[423] = out_r[23:8];
           result_i_ns[423] = out_i[23:8];
        end
        10'd87 : begin
           result_r_ns[935] = out_r[23:8];
           result_i_ns[935] = out_i[23:8];
        end
        10'd88 : begin
           result_r_ns[103] = out_r[23:8];
           result_i_ns[103] = out_i[23:8];
        end
        10'd89 : begin
           result_r_ns[615] = out_r[23:8];
           result_i_ns[615] = out_i[23:8];
        end
        10'd90 : begin
           result_r_ns[359] = out_r[23:8];
           result_i_ns[359] = out_i[23:8];
        end
        10'd91 : begin
           result_r_ns[871] = out_r[23:8];
           result_i_ns[871] = out_i[23:8];
        end
        10'd92 : begin
           result_r_ns[231] = out_r[23:8];
           result_i_ns[231] = out_i[23:8];
        end
        10'd93 : begin
           result_r_ns[743] = out_r[23:8];
           result_i_ns[743] = out_i[23:8];
        end
        10'd94 : begin
           result_r_ns[487] = out_r[23:8];
           result_i_ns[487] = out_i[23:8];
        end
        10'd95 : begin
           result_r_ns[999] = out_r[23:8];
           result_i_ns[999] = out_i[23:8];
        end
        10'd96 : begin
           result_r_ns[23] = out_r[23:8];
           result_i_ns[23] = out_i[23:8];
        end
        10'd97 : begin
           result_r_ns[535] = out_r[23:8];
           result_i_ns[535] = out_i[23:8];
        end
        10'd98 : begin
           result_r_ns[279] = out_r[23:8];
           result_i_ns[279] = out_i[23:8];
        end
        10'd99 : begin
           result_r_ns[791] = out_r[23:8];
           result_i_ns[791] = out_i[23:8];
        end
        10'd100 : begin
           result_r_ns[151] = out_r[23:8];
           result_i_ns[151] = out_i[23:8];
        end
        10'd101 : begin
           result_r_ns[663] = out_r[23:8];
           result_i_ns[663] = out_i[23:8];
        end
        10'd102 : begin
           result_r_ns[407] = out_r[23:8];
           result_i_ns[407] = out_i[23:8];
        end
        10'd103 : begin
           result_r_ns[919] = out_r[23:8];
           result_i_ns[919] = out_i[23:8];
        end
        10'd104 : begin
           result_r_ns[87] = out_r[23:8];
           result_i_ns[87] = out_i[23:8];
        end
        10'd105 : begin
           result_r_ns[599] = out_r[23:8];
           result_i_ns[599] = out_i[23:8];
        end
        10'd106 : begin
           result_r_ns[343] = out_r[23:8];
           result_i_ns[343] = out_i[23:8];
        end
        10'd107 : begin
           result_r_ns[855] = out_r[23:8];
           result_i_ns[855] = out_i[23:8];
        end
        10'd108 : begin
           result_r_ns[215] = out_r[23:8];
           result_i_ns[215] = out_i[23:8];
        end
        10'd109 : begin
           result_r_ns[727] = out_r[23:8];
           result_i_ns[727] = out_i[23:8];
        end
        10'd110 : begin
           result_r_ns[471] = out_r[23:8];
           result_i_ns[471] = out_i[23:8];
        end
        10'd111 : begin
           result_r_ns[983] = out_r[23:8];
           result_i_ns[983] = out_i[23:8];
        end
        10'd112 : begin
           result_r_ns[55] = out_r[23:8];
           result_i_ns[55] = out_i[23:8];
        end
        10'd113 : begin
           result_r_ns[567] = out_r[23:8];
           result_i_ns[567] = out_i[23:8];
        end
        10'd114 : begin
           result_r_ns[311] = out_r[23:8];
           result_i_ns[311] = out_i[23:8];
        end
        10'd115 : begin
           result_r_ns[823] = out_r[23:8];
           result_i_ns[823] = out_i[23:8];
        end
        10'd116 : begin
           result_r_ns[183] = out_r[23:8];
           result_i_ns[183] = out_i[23:8];
        end
        10'd117 : begin
           result_r_ns[695] = out_r[23:8];
           result_i_ns[695] = out_i[23:8];
        end
        10'd118 : begin
           result_r_ns[439] = out_r[23:8];
           result_i_ns[439] = out_i[23:8];
        end
        10'd119 : begin
           result_r_ns[951] = out_r[23:8];
           result_i_ns[951] = out_i[23:8];
        end
        10'd120 : begin
           result_r_ns[119] = out_r[23:8];
           result_i_ns[119] = out_i[23:8];
        end
        10'd121 : begin
           result_r_ns[631] = out_r[23:8];
           result_i_ns[631] = out_i[23:8];
        end
        10'd122 : begin
           result_r_ns[375] = out_r[23:8];
           result_i_ns[375] = out_i[23:8];
        end
        10'd123 : begin
           result_r_ns[887] = out_r[23:8];
           result_i_ns[887] = out_i[23:8];
        end
        10'd124 : begin
           result_r_ns[247] = out_r[23:8];
           result_i_ns[247] = out_i[23:8];
        end
        10'd125 : begin
           result_r_ns[759] = out_r[23:8];
           result_i_ns[759] = out_i[23:8];
        end
        10'd126 : begin
           result_r_ns[503] = out_r[23:8];
           result_i_ns[503] = out_i[23:8];
        end
        10'd127 : begin
           result_r_ns[1015] = out_r[23:8];
           result_i_ns[1015] = out_i[23:8];
        end
        10'd128 : begin
           result_r_ns[3] = out_r[23:8];
           result_i_ns[3] = out_i[23:8];
        end
        10'd129 : begin
           result_r_ns[515] = out_r[23:8];
           result_i_ns[515] = out_i[23:8];
        end
        10'd130 : begin
           result_r_ns[259] = out_r[23:8];
           result_i_ns[259] = out_i[23:8];
        end
        10'd131 : begin
           result_r_ns[771] = out_r[23:8];
           result_i_ns[771] = out_i[23:8];
        end
        10'd132 : begin
           result_r_ns[131] = out_r[23:8];
           result_i_ns[131] = out_i[23:8];
        end
        10'd133 : begin
           result_r_ns[643] = out_r[23:8];
           result_i_ns[643] = out_i[23:8];
        end
        10'd134 : begin
           result_r_ns[387] = out_r[23:8];
           result_i_ns[387] = out_i[23:8];
        end
        10'd135 : begin
           result_r_ns[899] = out_r[23:8];
           result_i_ns[899] = out_i[23:8];
        end
        10'd136 : begin
           result_r_ns[67] = out_r[23:8];
           result_i_ns[67] = out_i[23:8];
        end
        10'd137 : begin
           result_r_ns[579] = out_r[23:8];
           result_i_ns[579] = out_i[23:8];
        end
        10'd138 : begin
           result_r_ns[323] = out_r[23:8];
           result_i_ns[323] = out_i[23:8];
        end
        10'd139 : begin
           result_r_ns[835] = out_r[23:8];
           result_i_ns[835] = out_i[23:8];
        end
        10'd140 : begin
           result_r_ns[195] = out_r[23:8];
           result_i_ns[195] = out_i[23:8];
        end
        10'd141 : begin
           result_r_ns[707] = out_r[23:8];
           result_i_ns[707] = out_i[23:8];
        end
        10'd142 : begin
           result_r_ns[451] = out_r[23:8];
           result_i_ns[451] = out_i[23:8];
        end
        10'd143 : begin
           result_r_ns[963] = out_r[23:8];
           result_i_ns[963] = out_i[23:8];
        end
        10'd144 : begin
           result_r_ns[35] = out_r[23:8];
           result_i_ns[35] = out_i[23:8];
        end
        10'd145 : begin
           result_r_ns[547] = out_r[23:8];
           result_i_ns[547] = out_i[23:8];
        end
        10'd146 : begin
           result_r_ns[291] = out_r[23:8];
           result_i_ns[291] = out_i[23:8];
        end
        10'd147 : begin
           result_r_ns[803] = out_r[23:8];
           result_i_ns[803] = out_i[23:8];
        end
        10'd148 : begin
           result_r_ns[163] = out_r[23:8];
           result_i_ns[163] = out_i[23:8];
        end
        10'd149 : begin
           result_r_ns[675] = out_r[23:8];
           result_i_ns[675] = out_i[23:8];
        end
        10'd150 : begin
           result_r_ns[419] = out_r[23:8];
           result_i_ns[419] = out_i[23:8];
        end
        10'd151 : begin
           result_r_ns[931] = out_r[23:8];
           result_i_ns[931] = out_i[23:8];
        end
        10'd152 : begin
           result_r_ns[99] = out_r[23:8];
           result_i_ns[99] = out_i[23:8];
        end
        10'd153 : begin
           result_r_ns[611] = out_r[23:8];
           result_i_ns[611] = out_i[23:8];
        end
        10'd154 : begin
           result_r_ns[355] = out_r[23:8];
           result_i_ns[355] = out_i[23:8];
        end
        10'd155 : begin
           result_r_ns[867] = out_r[23:8];
           result_i_ns[867] = out_i[23:8];
        end
        10'd156 : begin
           result_r_ns[227] = out_r[23:8];
           result_i_ns[227] = out_i[23:8];
        end
        10'd157 : begin
           result_r_ns[739] = out_r[23:8];
           result_i_ns[739] = out_i[23:8];
        end
        10'd158 : begin
           result_r_ns[483] = out_r[23:8];
           result_i_ns[483] = out_i[23:8];
        end
        10'd159 : begin
           result_r_ns[995] = out_r[23:8];
           result_i_ns[995] = out_i[23:8];
        end
        10'd160 : begin
           result_r_ns[19] = out_r[23:8];
           result_i_ns[19] = out_i[23:8];
        end
        10'd161 : begin
           result_r_ns[531] = out_r[23:8];
           result_i_ns[531] = out_i[23:8];
        end
        10'd162 : begin
           result_r_ns[275] = out_r[23:8];
           result_i_ns[275] = out_i[23:8];
        end
        10'd163 : begin
           result_r_ns[787] = out_r[23:8];
           result_i_ns[787] = out_i[23:8];
        end
        10'd164 : begin
           result_r_ns[147] = out_r[23:8];
           result_i_ns[147] = out_i[23:8];
        end
        10'd165 : begin
           result_r_ns[659] = out_r[23:8];
           result_i_ns[659] = out_i[23:8];
        end
        10'd166 : begin
           result_r_ns[403] = out_r[23:8];
           result_i_ns[403] = out_i[23:8];
        end
        10'd167 : begin
           result_r_ns[915] = out_r[23:8];
           result_i_ns[915] = out_i[23:8];
        end
        10'd168 : begin
           result_r_ns[83] = out_r[23:8];
           result_i_ns[83] = out_i[23:8];
        end
        10'd169 : begin
           result_r_ns[595] = out_r[23:8];
           result_i_ns[595] = out_i[23:8];
        end
        10'd170 : begin
           result_r_ns[339] = out_r[23:8];
           result_i_ns[339] = out_i[23:8];
        end
        10'd171 : begin
           result_r_ns[851] = out_r[23:8];
           result_i_ns[851] = out_i[23:8];
        end
        10'd172 : begin
           result_r_ns[211] = out_r[23:8];
           result_i_ns[211] = out_i[23:8];
        end
        10'd173 : begin
           result_r_ns[723] = out_r[23:8];
           result_i_ns[723] = out_i[23:8];
        end
        10'd174 : begin
           result_r_ns[467] = out_r[23:8];
           result_i_ns[467] = out_i[23:8];
        end
        10'd175 : begin
           result_r_ns[979] = out_r[23:8];
           result_i_ns[979] = out_i[23:8];
        end
        10'd176 : begin
           result_r_ns[51] = out_r[23:8];
           result_i_ns[51] = out_i[23:8];
        end
        10'd177 : begin
           result_r_ns[563] = out_r[23:8];
           result_i_ns[563] = out_i[23:8];
        end
        10'd178 : begin
           result_r_ns[307] = out_r[23:8];
           result_i_ns[307] = out_i[23:8];
        end
        10'd179 : begin
           result_r_ns[819] = out_r[23:8];
           result_i_ns[819] = out_i[23:8];
        end
        10'd180 : begin
           result_r_ns[179] = out_r[23:8];
           result_i_ns[179] = out_i[23:8];
        end
        10'd181 : begin
           result_r_ns[691] = out_r[23:8];
           result_i_ns[691] = out_i[23:8];
        end
        10'd182 : begin
           result_r_ns[435] = out_r[23:8];
           result_i_ns[435] = out_i[23:8];
        end
        10'd183 : begin
           result_r_ns[947] = out_r[23:8];
           result_i_ns[947] = out_i[23:8];
        end
        10'd184 : begin
           result_r_ns[115] = out_r[23:8];
           result_i_ns[115] = out_i[23:8];
        end
        10'd185 : begin
           result_r_ns[627] = out_r[23:8];
           result_i_ns[627] = out_i[23:8];
        end
        10'd186 : begin
           result_r_ns[371] = out_r[23:8];
           result_i_ns[371] = out_i[23:8];
        end
        10'd187 : begin
           result_r_ns[883] = out_r[23:8];
           result_i_ns[883] = out_i[23:8];
        end
        10'd188 : begin
           result_r_ns[243] = out_r[23:8];
           result_i_ns[243] = out_i[23:8];
        end
        10'd189 : begin
           result_r_ns[755] = out_r[23:8];
           result_i_ns[755] = out_i[23:8];
        end
        10'd190 : begin
           result_r_ns[499] = out_r[23:8];
           result_i_ns[499] = out_i[23:8];
        end
        10'd191 : begin
           result_r_ns[1011] = out_r[23:8];
           result_i_ns[1011] = out_i[23:8];
        end
        10'd192 : begin
           result_r_ns[11] = out_r[23:8];
           result_i_ns[11] = out_i[23:8];
        end
        10'd193 : begin
           result_r_ns[523] = out_r[23:8];
           result_i_ns[523] = out_i[23:8];
        end
        10'd194 : begin
           result_r_ns[267] = out_r[23:8];
           result_i_ns[267] = out_i[23:8];
        end
        10'd195 : begin
           result_r_ns[779] = out_r[23:8];
           result_i_ns[779] = out_i[23:8];
        end
        10'd196 : begin
           result_r_ns[139] = out_r[23:8];
           result_i_ns[139] = out_i[23:8];
        end
        10'd197 : begin
           result_r_ns[651] = out_r[23:8];
           result_i_ns[651] = out_i[23:8];
        end
        10'd198 : begin
           result_r_ns[395] = out_r[23:8];
           result_i_ns[395] = out_i[23:8];
        end
        10'd199 : begin
           result_r_ns[907] = out_r[23:8];
           result_i_ns[907] = out_i[23:8];
        end
        10'd200 : begin
           result_r_ns[75] = out_r[23:8];
           result_i_ns[75] = out_i[23:8];
        end
        10'd201 : begin
           result_r_ns[587] = out_r[23:8];
           result_i_ns[587] = out_i[23:8];
        end
        10'd202 : begin
           result_r_ns[331] = out_r[23:8];
           result_i_ns[331] = out_i[23:8];
        end
        10'd203 : begin
           result_r_ns[843] = out_r[23:8];
           result_i_ns[843] = out_i[23:8];
        end
        10'd204 : begin
           result_r_ns[203] = out_r[23:8];
           result_i_ns[203] = out_i[23:8];
        end
        10'd205 : begin
           result_r_ns[715] = out_r[23:8];
           result_i_ns[715] = out_i[23:8];
        end
        10'd206 : begin
           result_r_ns[459] = out_r[23:8];
           result_i_ns[459] = out_i[23:8];
        end
        10'd207 : begin
           result_r_ns[971] = out_r[23:8];
           result_i_ns[971] = out_i[23:8];
        end
        10'd208 : begin
           result_r_ns[43] = out_r[23:8];
           result_i_ns[43] = out_i[23:8];
        end
        10'd209 : begin
           result_r_ns[555] = out_r[23:8];
           result_i_ns[555] = out_i[23:8];
        end
        10'd210 : begin
           result_r_ns[299] = out_r[23:8];
           result_i_ns[299] = out_i[23:8];
        end
        10'd211 : begin
           result_r_ns[811] = out_r[23:8];
           result_i_ns[811] = out_i[23:8];
        end
        10'd212 : begin
           result_r_ns[171] = out_r[23:8];
           result_i_ns[171] = out_i[23:8];
        end
        10'd213 : begin
           result_r_ns[683] = out_r[23:8];
           result_i_ns[683] = out_i[23:8];
        end
        10'd214 : begin
           result_r_ns[427] = out_r[23:8];
           result_i_ns[427] = out_i[23:8];
        end
        10'd215 : begin
           result_r_ns[939] = out_r[23:8];
           result_i_ns[939] = out_i[23:8];
        end
        10'd216 : begin
           result_r_ns[107] = out_r[23:8];
           result_i_ns[107] = out_i[23:8];
        end
        10'd217 : begin
           result_r_ns[619] = out_r[23:8];
           result_i_ns[619] = out_i[23:8];
        end
        10'd218 : begin
           result_r_ns[363] = out_r[23:8];
           result_i_ns[363] = out_i[23:8];
        end
        10'd219 : begin
           result_r_ns[875] = out_r[23:8];
           result_i_ns[875] = out_i[23:8];
        end
        10'd220 : begin
           result_r_ns[235] = out_r[23:8];
           result_i_ns[235] = out_i[23:8];
        end
        10'd221 : begin
           result_r_ns[747] = out_r[23:8];
           result_i_ns[747] = out_i[23:8];
        end
        10'd222 : begin
           result_r_ns[491] = out_r[23:8];
           result_i_ns[491] = out_i[23:8];
        end
        10'd223 : begin
           result_r_ns[1003] = out_r[23:8];
           result_i_ns[1003] = out_i[23:8];
        end
        10'd224 : begin
           result_r_ns[27] = out_r[23:8];
           result_i_ns[27] = out_i[23:8];
        end
        10'd225 : begin
           result_r_ns[539] = out_r[23:8];
           result_i_ns[539] = out_i[23:8];
        end
        10'd226 : begin
           result_r_ns[283] = out_r[23:8];
           result_i_ns[283] = out_i[23:8];
        end
        10'd227 : begin
           result_r_ns[795] = out_r[23:8];
           result_i_ns[795] = out_i[23:8];
        end
        10'd228 : begin
           result_r_ns[155] = out_r[23:8];
           result_i_ns[155] = out_i[23:8];
        end
        10'd229 : begin
           result_r_ns[667] = out_r[23:8];
           result_i_ns[667] = out_i[23:8];
        end
        10'd230 : begin
           result_r_ns[411] = out_r[23:8];
           result_i_ns[411] = out_i[23:8];
        end
        10'd231 : begin
           result_r_ns[923] = out_r[23:8];
           result_i_ns[923] = out_i[23:8];
        end
        10'd232 : begin
           result_r_ns[91] = out_r[23:8];
           result_i_ns[91] = out_i[23:8];
        end
        10'd233 : begin
           result_r_ns[603] = out_r[23:8];
           result_i_ns[603] = out_i[23:8];
        end
        10'd234 : begin
           result_r_ns[347] = out_r[23:8];
           result_i_ns[347] = out_i[23:8];
        end
        10'd235 : begin
           result_r_ns[859] = out_r[23:8];
           result_i_ns[859] = out_i[23:8];
        end
        10'd236 : begin
           result_r_ns[219] = out_r[23:8];
           result_i_ns[219] = out_i[23:8];
        end
        10'd237 : begin
           result_r_ns[731] = out_r[23:8];
           result_i_ns[731] = out_i[23:8];
        end
        10'd238 : begin
           result_r_ns[475] = out_r[23:8];
           result_i_ns[475] = out_i[23:8];
        end
        10'd239 : begin
           result_r_ns[987] = out_r[23:8];
           result_i_ns[987] = out_i[23:8];
        end
        10'd240 : begin
           result_r_ns[59] = out_r[23:8];
           result_i_ns[59] = out_i[23:8];
        end
        10'd241 : begin
           result_r_ns[571] = out_r[23:8];
           result_i_ns[571] = out_i[23:8];
        end
        10'd242 : begin
           result_r_ns[315] = out_r[23:8];
           result_i_ns[315] = out_i[23:8];
        end
        10'd243 : begin
           result_r_ns[827] = out_r[23:8];
           result_i_ns[827] = out_i[23:8];
        end
        10'd244 : begin
           result_r_ns[187] = out_r[23:8];
           result_i_ns[187] = out_i[23:8];
        end
        10'd245 : begin
           result_r_ns[699] = out_r[23:8];
           result_i_ns[699] = out_i[23:8];
        end
        10'd246 : begin
           result_r_ns[443] = out_r[23:8];
           result_i_ns[443] = out_i[23:8];
        end
        10'd247 : begin
           result_r_ns[955] = out_r[23:8];
           result_i_ns[955] = out_i[23:8];
        end
        10'd248 : begin
           result_r_ns[123] = out_r[23:8];
           result_i_ns[123] = out_i[23:8];
        end
        10'd249 : begin
           result_r_ns[635] = out_r[23:8];
           result_i_ns[635] = out_i[23:8];
        end
        10'd250 : begin
           result_r_ns[379] = out_r[23:8];
           result_i_ns[379] = out_i[23:8];
        end
        10'd251 : begin
           result_r_ns[891] = out_r[23:8];
           result_i_ns[891] = out_i[23:8];
        end
        10'd252 : begin
           result_r_ns[251] = out_r[23:8];
           result_i_ns[251] = out_i[23:8];
        end
        10'd253 : begin
           result_r_ns[763] = out_r[23:8];
           result_i_ns[763] = out_i[23:8];
        end
        10'd254 : begin
           result_r_ns[507] = out_r[23:8];
           result_i_ns[507] = out_i[23:8];
        end
        10'd255 : begin
           result_r_ns[1019] = out_r[23:8];
           result_i_ns[1019] = out_i[23:8];
        end
        10'd256 : begin
           result_r_ns[1] = out_r[23:8];
           result_i_ns[1] = out_i[23:8];
        end
        10'd257 : begin
           result_r_ns[513] = out_r[23:8];
           result_i_ns[513] = out_i[23:8];
        end
        10'd258 : begin
           result_r_ns[257] = out_r[23:8];
           result_i_ns[257] = out_i[23:8];
        end
        10'd259 : begin
           result_r_ns[769] = out_r[23:8];
           result_i_ns[769] = out_i[23:8];
        end
        10'd260 : begin
           result_r_ns[129] = out_r[23:8];
           result_i_ns[129] = out_i[23:8];
        end
        10'd261 : begin
           result_r_ns[641] = out_r[23:8];
           result_i_ns[641] = out_i[23:8];
        end
        10'd262 : begin
           result_r_ns[385] = out_r[23:8];
           result_i_ns[385] = out_i[23:8];
        end
        10'd263 : begin
           result_r_ns[897] = out_r[23:8];
           result_i_ns[897] = out_i[23:8];
        end
        10'd264 : begin
           result_r_ns[65] = out_r[23:8];
           result_i_ns[65] = out_i[23:8];
        end
        10'd265 : begin
           result_r_ns[577] = out_r[23:8];
           result_i_ns[577] = out_i[23:8];
        end
        10'd266 : begin
           result_r_ns[321] = out_r[23:8];
           result_i_ns[321] = out_i[23:8];
        end
        10'd267 : begin
           result_r_ns[833] = out_r[23:8];
           result_i_ns[833] = out_i[23:8];
        end
        10'd268 : begin
           result_r_ns[193] = out_r[23:8];
           result_i_ns[193] = out_i[23:8];
        end
        10'd269 : begin
           result_r_ns[705] = out_r[23:8];
           result_i_ns[705] = out_i[23:8];
        end
        10'd270 : begin
           result_r_ns[449] = out_r[23:8];
           result_i_ns[449] = out_i[23:8];
        end
        10'd271 : begin
           result_r_ns[961] = out_r[23:8];
           result_i_ns[961] = out_i[23:8];
        end
        10'd272 : begin
           result_r_ns[33] = out_r[23:8];
           result_i_ns[33] = out_i[23:8];
        end
        10'd273 : begin
           result_r_ns[545] = out_r[23:8];
           result_i_ns[545] = out_i[23:8];
        end
        10'd274 : begin
           result_r_ns[289] = out_r[23:8];
           result_i_ns[289] = out_i[23:8];
        end
        10'd275 : begin
           result_r_ns[801] = out_r[23:8];
           result_i_ns[801] = out_i[23:8];
        end
        10'd276 : begin
           result_r_ns[161] = out_r[23:8];
           result_i_ns[161] = out_i[23:8];
        end
        10'd277 : begin
           result_r_ns[673] = out_r[23:8];
           result_i_ns[673] = out_i[23:8];
        end
        10'd278 : begin
           result_r_ns[417] = out_r[23:8];
           result_i_ns[417] = out_i[23:8];
        end
        10'd279 : begin
           result_r_ns[929] = out_r[23:8];
           result_i_ns[929] = out_i[23:8];
        end
        10'd280 : begin
           result_r_ns[97] = out_r[23:8];
           result_i_ns[97] = out_i[23:8];
        end
        10'd281 : begin
           result_r_ns[609] = out_r[23:8];
           result_i_ns[609] = out_i[23:8];
        end
        10'd282 : begin
           result_r_ns[353] = out_r[23:8];
           result_i_ns[353] = out_i[23:8];
        end
        10'd283 : begin
           result_r_ns[865] = out_r[23:8];
           result_i_ns[865] = out_i[23:8];
        end
        10'd284 : begin
           result_r_ns[225] = out_r[23:8];
           result_i_ns[225] = out_i[23:8];
        end
        10'd285 : begin
           result_r_ns[737] = out_r[23:8];
           result_i_ns[737] = out_i[23:8];
        end
        10'd286 : begin
           result_r_ns[481] = out_r[23:8];
           result_i_ns[481] = out_i[23:8];
        end
        10'd287 : begin
           result_r_ns[993] = out_r[23:8];
           result_i_ns[993] = out_i[23:8];
        end
        10'd288 : begin
           result_r_ns[17] = out_r[23:8];
           result_i_ns[17] = out_i[23:8];
        end
        10'd289 : begin
           result_r_ns[529] = out_r[23:8];
           result_i_ns[529] = out_i[23:8];
        end
        10'd290 : begin
           result_r_ns[273] = out_r[23:8];
           result_i_ns[273] = out_i[23:8];
        end
        10'd291 : begin
           result_r_ns[785] = out_r[23:8];
           result_i_ns[785] = out_i[23:8];
        end
        10'd292 : begin
           result_r_ns[145] = out_r[23:8];
           result_i_ns[145] = out_i[23:8];
        end
        10'd293 : begin
           result_r_ns[657] = out_r[23:8];
           result_i_ns[657] = out_i[23:8];
        end
        10'd294 : begin
           result_r_ns[401] = out_r[23:8];
           result_i_ns[401] = out_i[23:8];
        end
        10'd295 : begin
           result_r_ns[913] = out_r[23:8];
           result_i_ns[913] = out_i[23:8];
        end
        10'd296 : begin
           result_r_ns[81] = out_r[23:8];
           result_i_ns[81] = out_i[23:8];
        end
        10'd297 : begin
           result_r_ns[593] = out_r[23:8];
           result_i_ns[593] = out_i[23:8];
        end
        10'd298 : begin
           result_r_ns[337] = out_r[23:8];
           result_i_ns[337] = out_i[23:8];
        end
        10'd299 : begin
           result_r_ns[849] = out_r[23:8];
           result_i_ns[849] = out_i[23:8];
        end
        10'd300 : begin
           result_r_ns[209] = out_r[23:8];
           result_i_ns[209] = out_i[23:8];
        end
        10'd301 : begin
           result_r_ns[721] = out_r[23:8];
           result_i_ns[721] = out_i[23:8];
        end
        10'd302 : begin
           result_r_ns[465] = out_r[23:8];
           result_i_ns[465] = out_i[23:8];
        end
        10'd303 : begin
           result_r_ns[977] = out_r[23:8];
           result_i_ns[977] = out_i[23:8];
        end
        10'd304 : begin
           result_r_ns[49] = out_r[23:8];
           result_i_ns[49] = out_i[23:8];
        end
        10'd305 : begin
           result_r_ns[561] = out_r[23:8];
           result_i_ns[561] = out_i[23:8];
        end
        10'd306 : begin
           result_r_ns[305] = out_r[23:8];
           result_i_ns[305] = out_i[23:8];
        end
        10'd307 : begin
           result_r_ns[817] = out_r[23:8];
           result_i_ns[817] = out_i[23:8];
        end
        10'd308 : begin
           result_r_ns[177] = out_r[23:8];
           result_i_ns[177] = out_i[23:8];
        end
        10'd309 : begin
           result_r_ns[689] = out_r[23:8];
           result_i_ns[689] = out_i[23:8];
        end
        10'd310 : begin
           result_r_ns[433] = out_r[23:8];
           result_i_ns[433] = out_i[23:8];
        end
        10'd311 : begin
           result_r_ns[945] = out_r[23:8];
           result_i_ns[945] = out_i[23:8];
        end
        10'd312 : begin
           result_r_ns[113] = out_r[23:8];
           result_i_ns[113] = out_i[23:8];
        end
        10'd313 : begin
           result_r_ns[625] = out_r[23:8];
           result_i_ns[625] = out_i[23:8];
        end
        10'd314 : begin
           result_r_ns[369] = out_r[23:8];
           result_i_ns[369] = out_i[23:8];
        end
        10'd315 : begin
           result_r_ns[881] = out_r[23:8];
           result_i_ns[881] = out_i[23:8];
        end
        10'd316 : begin
           result_r_ns[241] = out_r[23:8];
           result_i_ns[241] = out_i[23:8];
        end
        10'd317 : begin
           result_r_ns[753] = out_r[23:8];
           result_i_ns[753] = out_i[23:8];
        end
        10'd318 : begin
           result_r_ns[497] = out_r[23:8];
           result_i_ns[497] = out_i[23:8];
        end
        10'd319 : begin
           result_r_ns[1009] = out_r[23:8];
           result_i_ns[1009] = out_i[23:8];
        end
        10'd320 : begin
           result_r_ns[9] = out_r[23:8];
           result_i_ns[9] = out_i[23:8];
        end
        10'd321 : begin
           result_r_ns[521] = out_r[23:8];
           result_i_ns[521] = out_i[23:8];
        end
        10'd322 : begin
           result_r_ns[265] = out_r[23:8];
           result_i_ns[265] = out_i[23:8];
        end
        10'd323 : begin
           result_r_ns[777] = out_r[23:8];
           result_i_ns[777] = out_i[23:8];
        end
        10'd324 : begin
           result_r_ns[137] = out_r[23:8];
           result_i_ns[137] = out_i[23:8];
        end
        10'd325 : begin
           result_r_ns[649] = out_r[23:8];
           result_i_ns[649] = out_i[23:8];
        end
        10'd326 : begin
           result_r_ns[393] = out_r[23:8];
           result_i_ns[393] = out_i[23:8];
        end
        10'd327 : begin
           result_r_ns[905] = out_r[23:8];
           result_i_ns[905] = out_i[23:8];
        end
        10'd328 : begin
           result_r_ns[73] = out_r[23:8];
           result_i_ns[73] = out_i[23:8];
        end
        10'd329 : begin
           result_r_ns[585] = out_r[23:8];
           result_i_ns[585] = out_i[23:8];
        end
        10'd330 : begin
           result_r_ns[329] = out_r[23:8];
           result_i_ns[329] = out_i[23:8];
        end
        10'd331 : begin
           result_r_ns[841] = out_r[23:8];
           result_i_ns[841] = out_i[23:8];
        end
        10'd332 : begin
           result_r_ns[201] = out_r[23:8];
           result_i_ns[201] = out_i[23:8];
        end
        10'd333 : begin
           result_r_ns[713] = out_r[23:8];
           result_i_ns[713] = out_i[23:8];
        end
        10'd334 : begin
           result_r_ns[457] = out_r[23:8];
           result_i_ns[457] = out_i[23:8];
        end
        10'd335 : begin
           result_r_ns[969] = out_r[23:8];
           result_i_ns[969] = out_i[23:8];
        end
        10'd336 : begin
           result_r_ns[41] = out_r[23:8];
           result_i_ns[41] = out_i[23:8];
        end
        10'd337 : begin
           result_r_ns[553] = out_r[23:8];
           result_i_ns[553] = out_i[23:8];
        end
        10'd338 : begin
           result_r_ns[297] = out_r[23:8];
           result_i_ns[297] = out_i[23:8];
        end
        10'd339 : begin
           result_r_ns[809] = out_r[23:8];
           result_i_ns[809] = out_i[23:8];
        end
        10'd340 : begin
           result_r_ns[169] = out_r[23:8];
           result_i_ns[169] = out_i[23:8];
        end
        10'd341 : begin
           result_r_ns[681] = out_r[23:8];
           result_i_ns[681] = out_i[23:8];
        end
        10'd342 : begin
           result_r_ns[425] = out_r[23:8];
           result_i_ns[425] = out_i[23:8];
        end
        10'd343 : begin
           result_r_ns[937] = out_r[23:8];
           result_i_ns[937] = out_i[23:8];
        end
        10'd344 : begin
           result_r_ns[105] = out_r[23:8];
           result_i_ns[105] = out_i[23:8];
        end
        10'd345 : begin
           result_r_ns[617] = out_r[23:8];
           result_i_ns[617] = out_i[23:8];
        end
        10'd346 : begin
           result_r_ns[361] = out_r[23:8];
           result_i_ns[361] = out_i[23:8];
        end
        10'd347 : begin
           result_r_ns[873] = out_r[23:8];
           result_i_ns[873] = out_i[23:8];
        end
        10'd348 : begin
           result_r_ns[233] = out_r[23:8];
           result_i_ns[233] = out_i[23:8];
        end
        10'd349 : begin
           result_r_ns[745] = out_r[23:8];
           result_i_ns[745] = out_i[23:8];
        end
        10'd350 : begin
           result_r_ns[489] = out_r[23:8];
           result_i_ns[489] = out_i[23:8];
        end
        10'd351 : begin
           result_r_ns[1001] = out_r[23:8];
           result_i_ns[1001] = out_i[23:8];
        end
        10'd352 : begin
           result_r_ns[25] = out_r[23:8];
           result_i_ns[25] = out_i[23:8];
        end
        10'd353 : begin
           result_r_ns[537] = out_r[23:8];
           result_i_ns[537] = out_i[23:8];
        end
        10'd354 : begin
           result_r_ns[281] = out_r[23:8];
           result_i_ns[281] = out_i[23:8];
        end
        10'd355 : begin
           result_r_ns[793] = out_r[23:8];
           result_i_ns[793] = out_i[23:8];
        end
        10'd356 : begin
           result_r_ns[153] = out_r[23:8];
           result_i_ns[153] = out_i[23:8];
        end
        10'd357 : begin
           result_r_ns[665] = out_r[23:8];
           result_i_ns[665] = out_i[23:8];
        end
        10'd358 : begin
           result_r_ns[409] = out_r[23:8];
           result_i_ns[409] = out_i[23:8];
        end
        10'd359 : begin
           result_r_ns[921] = out_r[23:8];
           result_i_ns[921] = out_i[23:8];
        end
        10'd360 : begin
           result_r_ns[89] = out_r[23:8];
           result_i_ns[89] = out_i[23:8];
        end
        10'd361 : begin
           result_r_ns[601] = out_r[23:8];
           result_i_ns[601] = out_i[23:8];
        end
        10'd362 : begin
           result_r_ns[345] = out_r[23:8];
           result_i_ns[345] = out_i[23:8];
        end
        10'd363 : begin
           result_r_ns[857] = out_r[23:8];
           result_i_ns[857] = out_i[23:8];
        end
        10'd364 : begin
           result_r_ns[217] = out_r[23:8];
           result_i_ns[217] = out_i[23:8];
        end
        10'd365 : begin
           result_r_ns[729] = out_r[23:8];
           result_i_ns[729] = out_i[23:8];
        end
        10'd366 : begin
           result_r_ns[473] = out_r[23:8];
           result_i_ns[473] = out_i[23:8];
        end
        10'd367 : begin
           result_r_ns[985] = out_r[23:8];
           result_i_ns[985] = out_i[23:8];
        end
        10'd368 : begin
           result_r_ns[57] = out_r[23:8];
           result_i_ns[57] = out_i[23:8];
        end
        10'd369 : begin
           result_r_ns[569] = out_r[23:8];
           result_i_ns[569] = out_i[23:8];
        end
        10'd370 : begin
           result_r_ns[313] = out_r[23:8];
           result_i_ns[313] = out_i[23:8];
        end
        10'd371 : begin
           result_r_ns[825] = out_r[23:8];
           result_i_ns[825] = out_i[23:8];
        end
        10'd372 : begin
           result_r_ns[185] = out_r[23:8];
           result_i_ns[185] = out_i[23:8];
        end
        10'd373 : begin
           result_r_ns[697] = out_r[23:8];
           result_i_ns[697] = out_i[23:8];
        end
        10'd374 : begin
           result_r_ns[441] = out_r[23:8];
           result_i_ns[441] = out_i[23:8];
        end
        10'd375 : begin
           result_r_ns[953] = out_r[23:8];
           result_i_ns[953] = out_i[23:8];
        end
        10'd376 : begin
           result_r_ns[121] = out_r[23:8];
           result_i_ns[121] = out_i[23:8];
        end
        10'd377 : begin
           result_r_ns[633] = out_r[23:8];
           result_i_ns[633] = out_i[23:8];
        end
        10'd378 : begin
           result_r_ns[377] = out_r[23:8];
           result_i_ns[377] = out_i[23:8];
        end
        10'd379 : begin
           result_r_ns[889] = out_r[23:8];
           result_i_ns[889] = out_i[23:8];
        end
        10'd380 : begin
           result_r_ns[249] = out_r[23:8];
           result_i_ns[249] = out_i[23:8];
        end
        10'd381 : begin
           result_r_ns[761] = out_r[23:8];
           result_i_ns[761] = out_i[23:8];
        end
        10'd382 : begin
           result_r_ns[505] = out_r[23:8];
           result_i_ns[505] = out_i[23:8];
        end
        10'd383 : begin
           result_r_ns[1017] = out_r[23:8];
           result_i_ns[1017] = out_i[23:8];
        end
        10'd384 : begin
           result_r_ns[5] = out_r[23:8];
           result_i_ns[5] = out_i[23:8];
        end
        10'd385 : begin
           result_r_ns[517] = out_r[23:8];
           result_i_ns[517] = out_i[23:8];
        end
        10'd386 : begin
           result_r_ns[261] = out_r[23:8];
           result_i_ns[261] = out_i[23:8];
        end
        10'd387 : begin
           result_r_ns[773] = out_r[23:8];
           result_i_ns[773] = out_i[23:8];
        end
        10'd388 : begin
           result_r_ns[133] = out_r[23:8];
           result_i_ns[133] = out_i[23:8];
        end
        10'd389 : begin
           result_r_ns[645] = out_r[23:8];
           result_i_ns[645] = out_i[23:8];
        end
        10'd390 : begin
           result_r_ns[389] = out_r[23:8];
           result_i_ns[389] = out_i[23:8];
        end
        10'd391 : begin
           result_r_ns[901] = out_r[23:8];
           result_i_ns[901] = out_i[23:8];
        end
        10'd392 : begin
           result_r_ns[69] = out_r[23:8];
           result_i_ns[69] = out_i[23:8];
        end
        10'd393 : begin
           result_r_ns[581] = out_r[23:8];
           result_i_ns[581] = out_i[23:8];
        end
        10'd394 : begin
           result_r_ns[325] = out_r[23:8];
           result_i_ns[325] = out_i[23:8];
        end
        10'd395 : begin
           result_r_ns[837] = out_r[23:8];
           result_i_ns[837] = out_i[23:8];
        end
        10'd396 : begin
           result_r_ns[197] = out_r[23:8];
           result_i_ns[197] = out_i[23:8];
        end
        10'd397 : begin
           result_r_ns[709] = out_r[23:8];
           result_i_ns[709] = out_i[23:8];
        end
        10'd398 : begin
           result_r_ns[453] = out_r[23:8];
           result_i_ns[453] = out_i[23:8];
        end
        10'd399 : begin
           result_r_ns[965] = out_r[23:8];
           result_i_ns[965] = out_i[23:8];
        end
        10'd400 : begin
           result_r_ns[37] = out_r[23:8];
           result_i_ns[37] = out_i[23:8];
        end
        10'd401 : begin
           result_r_ns[549] = out_r[23:8];
           result_i_ns[549] = out_i[23:8];
        end
        10'd402 : begin
           result_r_ns[293] = out_r[23:8];
           result_i_ns[293] = out_i[23:8];
        end
        10'd403 : begin
           result_r_ns[805] = out_r[23:8];
           result_i_ns[805] = out_i[23:8];
        end
        10'd404 : begin
           result_r_ns[165] = out_r[23:8];
           result_i_ns[165] = out_i[23:8];
        end
        10'd405 : begin
           result_r_ns[677] = out_r[23:8];
           result_i_ns[677] = out_i[23:8];
        end
        10'd406 : begin
           result_r_ns[421] = out_r[23:8];
           result_i_ns[421] = out_i[23:8];
        end
        10'd407 : begin
           result_r_ns[933] = out_r[23:8];
           result_i_ns[933] = out_i[23:8];
        end
        10'd408 : begin
           result_r_ns[101] = out_r[23:8];
           result_i_ns[101] = out_i[23:8];
        end
        10'd409 : begin
           result_r_ns[613] = out_r[23:8];
           result_i_ns[613] = out_i[23:8];
        end
        10'd410 : begin
           result_r_ns[357] = out_r[23:8];
           result_i_ns[357] = out_i[23:8];
        end
        10'd411 : begin
           result_r_ns[869] = out_r[23:8];
           result_i_ns[869] = out_i[23:8];
        end
        10'd412 : begin
           result_r_ns[229] = out_r[23:8];
           result_i_ns[229] = out_i[23:8];
        end
        10'd413 : begin
           result_r_ns[741] = out_r[23:8];
           result_i_ns[741] = out_i[23:8];
        end
        10'd414 : begin
           result_r_ns[485] = out_r[23:8];
           result_i_ns[485] = out_i[23:8];
        end
        10'd415 : begin
           result_r_ns[997] = out_r[23:8];
           result_i_ns[997] = out_i[23:8];
        end
        10'd416 : begin
           result_r_ns[21] = out_r[23:8];
           result_i_ns[21] = out_i[23:8];
        end
        10'd417 : begin
           result_r_ns[533] = out_r[23:8];
           result_i_ns[533] = out_i[23:8];
        end
        10'd418 : begin
           result_r_ns[277] = out_r[23:8];
           result_i_ns[277] = out_i[23:8];
        end
        10'd419 : begin
           result_r_ns[789] = out_r[23:8];
           result_i_ns[789] = out_i[23:8];
        end
        10'd420 : begin
           result_r_ns[149] = out_r[23:8];
           result_i_ns[149] = out_i[23:8];
        end
        10'd421 : begin
           result_r_ns[661] = out_r[23:8];
           result_i_ns[661] = out_i[23:8];
        end
        10'd422 : begin
           result_r_ns[405] = out_r[23:8];
           result_i_ns[405] = out_i[23:8];
        end
        10'd423 : begin
           result_r_ns[917] = out_r[23:8];
           result_i_ns[917] = out_i[23:8];
        end
        10'd424 : begin
           result_r_ns[85] = out_r[23:8];
           result_i_ns[85] = out_i[23:8];
        end
        10'd425 : begin
           result_r_ns[597] = out_r[23:8];
           result_i_ns[597] = out_i[23:8];
        end
        10'd426 : begin
           result_r_ns[341] = out_r[23:8];
           result_i_ns[341] = out_i[23:8];
        end
        10'd427 : begin
           result_r_ns[853] = out_r[23:8];
           result_i_ns[853] = out_i[23:8];
        end
        10'd428 : begin
           result_r_ns[213] = out_r[23:8];
           result_i_ns[213] = out_i[23:8];
        end
        10'd429 : begin
           result_r_ns[725] = out_r[23:8];
           result_i_ns[725] = out_i[23:8];
        end
        10'd430 : begin
           result_r_ns[469] = out_r[23:8];
           result_i_ns[469] = out_i[23:8];
        end
        10'd431 : begin
           result_r_ns[981] = out_r[23:8];
           result_i_ns[981] = out_i[23:8];
        end
        10'd432 : begin
           result_r_ns[53] = out_r[23:8];
           result_i_ns[53] = out_i[23:8];
        end
        10'd433 : begin
           result_r_ns[565] = out_r[23:8];
           result_i_ns[565] = out_i[23:8];
        end
        10'd434 : begin
           result_r_ns[309] = out_r[23:8];
           result_i_ns[309] = out_i[23:8];
        end
        10'd435 : begin
           result_r_ns[821] = out_r[23:8];
           result_i_ns[821] = out_i[23:8];
        end
        10'd436 : begin
           result_r_ns[181] = out_r[23:8];
           result_i_ns[181] = out_i[23:8];
        end
        10'd437 : begin
           result_r_ns[693] = out_r[23:8];
           result_i_ns[693] = out_i[23:8];
        end
        10'd438 : begin
           result_r_ns[437] = out_r[23:8];
           result_i_ns[437] = out_i[23:8];
        end
        10'd439 : begin
           result_r_ns[949] = out_r[23:8];
           result_i_ns[949] = out_i[23:8];
        end
        10'd440 : begin
           result_r_ns[117] = out_r[23:8];
           result_i_ns[117] = out_i[23:8];
        end
        10'd441 : begin
           result_r_ns[629] = out_r[23:8];
           result_i_ns[629] = out_i[23:8];
        end
        10'd442 : begin
           result_r_ns[373] = out_r[23:8];
           result_i_ns[373] = out_i[23:8];
        end
        10'd443 : begin
           result_r_ns[885] = out_r[23:8];
           result_i_ns[885] = out_i[23:8];
        end
        10'd444 : begin
           result_r_ns[245] = out_r[23:8];
           result_i_ns[245] = out_i[23:8];
        end
        10'd445 : begin
           result_r_ns[757] = out_r[23:8];
           result_i_ns[757] = out_i[23:8];
        end
        10'd446 : begin
           result_r_ns[501] = out_r[23:8];
           result_i_ns[501] = out_i[23:8];
        end
        10'd447 : begin
           result_r_ns[1013] = out_r[23:8];
           result_i_ns[1013] = out_i[23:8];
        end
        10'd448 : begin
           result_r_ns[13] = out_r[23:8];
           result_i_ns[13] = out_i[23:8];
        end
        10'd449 : begin
           result_r_ns[525] = out_r[23:8];
           result_i_ns[525] = out_i[23:8];
        end
        10'd450 : begin
           result_r_ns[269] = out_r[23:8];
           result_i_ns[269] = out_i[23:8];
        end
        10'd451 : begin
           result_r_ns[781] = out_r[23:8];
           result_i_ns[781] = out_i[23:8];
        end
        10'd452 : begin
           result_r_ns[141] = out_r[23:8];
           result_i_ns[141] = out_i[23:8];
        end
        10'd453 : begin
           result_r_ns[653] = out_r[23:8];
           result_i_ns[653] = out_i[23:8];
        end
        10'd454 : begin
           result_r_ns[397] = out_r[23:8];
           result_i_ns[397] = out_i[23:8];
        end
        10'd455 : begin
           result_r_ns[909] = out_r[23:8];
           result_i_ns[909] = out_i[23:8];
        end
        10'd456 : begin
           result_r_ns[77] = out_r[23:8];
           result_i_ns[77] = out_i[23:8];
        end
        10'd457 : begin
           result_r_ns[589] = out_r[23:8];
           result_i_ns[589] = out_i[23:8];
        end
        10'd458 : begin
           result_r_ns[333] = out_r[23:8];
           result_i_ns[333] = out_i[23:8];
        end
        10'd459 : begin
           result_r_ns[845] = out_r[23:8];
           result_i_ns[845] = out_i[23:8];
        end
        10'd460 : begin
           result_r_ns[205] = out_r[23:8];
           result_i_ns[205] = out_i[23:8];
        end
        10'd461 : begin
           result_r_ns[717] = out_r[23:8];
           result_i_ns[717] = out_i[23:8];
        end
        10'd462 : begin
           result_r_ns[461] = out_r[23:8];
           result_i_ns[461] = out_i[23:8];
        end
        10'd463 : begin
           result_r_ns[973] = out_r[23:8];
           result_i_ns[973] = out_i[23:8];
        end
        10'd464 : begin
           result_r_ns[45] = out_r[23:8];
           result_i_ns[45] = out_i[23:8];
        end
        10'd465 : begin
           result_r_ns[557] = out_r[23:8];
           result_i_ns[557] = out_i[23:8];
        end
        10'd466 : begin
           result_r_ns[301] = out_r[23:8];
           result_i_ns[301] = out_i[23:8];
        end
        10'd467 : begin
           result_r_ns[813] = out_r[23:8];
           result_i_ns[813] = out_i[23:8];
        end
        10'd468 : begin
           result_r_ns[173] = out_r[23:8];
           result_i_ns[173] = out_i[23:8];
        end
        10'd469 : begin
           result_r_ns[685] = out_r[23:8];
           result_i_ns[685] = out_i[23:8];
        end
        10'd470 : begin
           result_r_ns[429] = out_r[23:8];
           result_i_ns[429] = out_i[23:8];
        end
        10'd471 : begin
           result_r_ns[941] = out_r[23:8];
           result_i_ns[941] = out_i[23:8];
        end
        10'd472 : begin
           result_r_ns[109] = out_r[23:8];
           result_i_ns[109] = out_i[23:8];
        end
        10'd473 : begin
           result_r_ns[621] = out_r[23:8];
           result_i_ns[621] = out_i[23:8];
        end
        10'd474 : begin
           result_r_ns[365] = out_r[23:8];
           result_i_ns[365] = out_i[23:8];
        end
        10'd475 : begin
           result_r_ns[877] = out_r[23:8];
           result_i_ns[877] = out_i[23:8];
        end
        10'd476 : begin
           result_r_ns[237] = out_r[23:8];
           result_i_ns[237] = out_i[23:8];
        end
        10'd477 : begin
           result_r_ns[749] = out_r[23:8];
           result_i_ns[749] = out_i[23:8];
        end
        10'd478 : begin
           result_r_ns[493] = out_r[23:8];
           result_i_ns[493] = out_i[23:8];
        end
        10'd479 : begin
           result_r_ns[1005] = out_r[23:8];
           result_i_ns[1005] = out_i[23:8];
        end
        10'd480 : begin
           result_r_ns[29] = out_r[23:8];
           result_i_ns[29] = out_i[23:8];
        end
        10'd481 : begin
           result_r_ns[541] = out_r[23:8];
           result_i_ns[541] = out_i[23:8];
        end
        10'd482 : begin
           result_r_ns[285] = out_r[23:8];
           result_i_ns[285] = out_i[23:8];
        end
        10'd483 : begin
           result_r_ns[797] = out_r[23:8];
           result_i_ns[797] = out_i[23:8];
        end
        10'd484 : begin
           result_r_ns[157] = out_r[23:8];
           result_i_ns[157] = out_i[23:8];
        end
        10'd485 : begin
           result_r_ns[669] = out_r[23:8];
           result_i_ns[669] = out_i[23:8];
        end
        10'd486 : begin
           result_r_ns[413] = out_r[23:8];
           result_i_ns[413] = out_i[23:8];
        end
        10'd487 : begin
           result_r_ns[925] = out_r[23:8];
           result_i_ns[925] = out_i[23:8];
        end
        10'd488 : begin
           result_r_ns[93] = out_r[23:8];
           result_i_ns[93] = out_i[23:8];
        end
        10'd489 : begin
           result_r_ns[605] = out_r[23:8];
           result_i_ns[605] = out_i[23:8];
        end
        10'd490 : begin
           result_r_ns[349] = out_r[23:8];
           result_i_ns[349] = out_i[23:8];
        end
        10'd491 : begin
           result_r_ns[861] = out_r[23:8];
           result_i_ns[861] = out_i[23:8];
        end
        10'd492 : begin
           result_r_ns[221] = out_r[23:8];
           result_i_ns[221] = out_i[23:8];
        end
        10'd493 : begin
           result_r_ns[733] = out_r[23:8];
           result_i_ns[733] = out_i[23:8];
        end
        10'd494 : begin
           result_r_ns[477] = out_r[23:8];
           result_i_ns[477] = out_i[23:8];
        end
        10'd495 : begin
           result_r_ns[989] = out_r[23:8];
           result_i_ns[989] = out_i[23:8];
        end
        10'd496 : begin
           result_r_ns[61] = out_r[23:8];
           result_i_ns[61] = out_i[23:8];
        end
        10'd497 : begin
           result_r_ns[573] = out_r[23:8];
           result_i_ns[573] = out_i[23:8];
        end
        10'd498 : begin
           result_r_ns[317] = out_r[23:8];
           result_i_ns[317] = out_i[23:8];
        end
        10'd499 : begin
           result_r_ns[829] = out_r[23:8];
           result_i_ns[829] = out_i[23:8];
        end
        10'd500 : begin
           result_r_ns[189] = out_r[23:8];
           result_i_ns[189] = out_i[23:8];
        end
        10'd501 : begin
           result_r_ns[701] = out_r[23:8];
           result_i_ns[701] = out_i[23:8];
        end
        10'd502 : begin
           result_r_ns[445] = out_r[23:8];
           result_i_ns[445] = out_i[23:8];
        end
        10'd503 : begin
           result_r_ns[957] = out_r[23:8];
           result_i_ns[957] = out_i[23:8];
        end
        10'd504 : begin
           result_r_ns[125] = out_r[23:8];
           result_i_ns[125] = out_i[23:8];
        end
        10'd505 : begin
           result_r_ns[637] = out_r[23:8];
           result_i_ns[637] = out_i[23:8];
        end
        10'd506 : begin
           result_r_ns[381] = out_r[23:8];
           result_i_ns[381] = out_i[23:8];
        end
        10'd507 : begin
           result_r_ns[893] = out_r[23:8];
           result_i_ns[893] = out_i[23:8];
        end
        10'd508 : begin
           result_r_ns[253] = out_r[23:8];
           result_i_ns[253] = out_i[23:8];
        end
        10'd509 : begin
           result_r_ns[765] = out_r[23:8];
           result_i_ns[765] = out_i[23:8];
        end
        10'd510 : begin
           result_r_ns[509] = out_r[23:8];
           result_i_ns[509] = out_i[23:8];
        end
        10'd511 : begin
           result_r_ns[1021] = out_r[23:8];
           result_i_ns[1021] = out_i[23:8];
        end
        10'd512 : begin
           result_r_ns[0] = out_r[23:8];
           result_i_ns[0] = out_i[23:8];
        end
        10'd513 : begin
           result_r_ns[512] = out_r[23:8];
           result_i_ns[512] = out_i[23:8];
        end
        10'd514 : begin
           result_r_ns[256] = out_r[23:8];
           result_i_ns[256] = out_i[23:8];
        end
        10'd515 : begin
           result_r_ns[768] = out_r[23:8];
           result_i_ns[768] = out_i[23:8];
        end
        10'd516 : begin
           result_r_ns[128] = out_r[23:8];
           result_i_ns[128] = out_i[23:8];
        end
        10'd517 : begin
           result_r_ns[640] = out_r[23:8];
           result_i_ns[640] = out_i[23:8];
        end
        10'd518 : begin
           result_r_ns[384] = out_r[23:8];
           result_i_ns[384] = out_i[23:8];
        end
        10'd519 : begin
           result_r_ns[896] = out_r[23:8];
           result_i_ns[896] = out_i[23:8];
        end
        10'd520 : begin
           result_r_ns[64] = out_r[23:8];
           result_i_ns[64] = out_i[23:8];
        end
        10'd521 : begin
           result_r_ns[576] = out_r[23:8];
           result_i_ns[576] = out_i[23:8];
        end
        10'd522 : begin
           result_r_ns[320] = out_r[23:8];
           result_i_ns[320] = out_i[23:8];
        end
        10'd523 : begin
           result_r_ns[832] = out_r[23:8];
           result_i_ns[832] = out_i[23:8];
        end
        10'd524 : begin
           result_r_ns[192] = out_r[23:8];
           result_i_ns[192] = out_i[23:8];
        end
        10'd525 : begin
           result_r_ns[704] = out_r[23:8];
           result_i_ns[704] = out_i[23:8];
        end
        10'd526 : begin
           result_r_ns[448] = out_r[23:8];
           result_i_ns[448] = out_i[23:8];
        end
        10'd527 : begin
           result_r_ns[960] = out_r[23:8];
           result_i_ns[960] = out_i[23:8];
        end
        10'd528 : begin
           result_r_ns[32] = out_r[23:8];
           result_i_ns[32] = out_i[23:8];
        end
        10'd529 : begin
           result_r_ns[544] = out_r[23:8];
           result_i_ns[544] = out_i[23:8];
        end
        10'd530 : begin
           result_r_ns[288] = out_r[23:8];
           result_i_ns[288] = out_i[23:8];
        end
        10'd531 : begin
           result_r_ns[800] = out_r[23:8];
           result_i_ns[800] = out_i[23:8];
        end
        10'd532 : begin
           result_r_ns[160] = out_r[23:8];
           result_i_ns[160] = out_i[23:8];
        end
        10'd533 : begin
           result_r_ns[672] = out_r[23:8];
           result_i_ns[672] = out_i[23:8];
        end
        10'd534 : begin
           result_r_ns[416] = out_r[23:8];
           result_i_ns[416] = out_i[23:8];
        end
        10'd535 : begin
           result_r_ns[928] = out_r[23:8];
           result_i_ns[928] = out_i[23:8];
        end
        10'd536 : begin
           result_r_ns[96] = out_r[23:8];
           result_i_ns[96] = out_i[23:8];
        end
        10'd537 : begin
           result_r_ns[608] = out_r[23:8];
           result_i_ns[608] = out_i[23:8];
        end
        10'd538 : begin
           result_r_ns[352] = out_r[23:8];
           result_i_ns[352] = out_i[23:8];
        end
        10'd539 : begin
           result_r_ns[864] = out_r[23:8];
           result_i_ns[864] = out_i[23:8];
        end
        10'd540 : begin
           result_r_ns[224] = out_r[23:8];
           result_i_ns[224] = out_i[23:8];
        end
        10'd541 : begin
           result_r_ns[736] = out_r[23:8];
           result_i_ns[736] = out_i[23:8];
        end
        10'd542 : begin
           result_r_ns[480] = out_r[23:8];
           result_i_ns[480] = out_i[23:8];
        end
        10'd543 : begin
           result_r_ns[992] = out_r[23:8];
           result_i_ns[992] = out_i[23:8];
        end
        10'd544 : begin
           result_r_ns[16] = out_r[23:8];
           result_i_ns[16] = out_i[23:8];
        end
        10'd545 : begin
           result_r_ns[528] = out_r[23:8];
           result_i_ns[528] = out_i[23:8];
        end
        10'd546 : begin
           result_r_ns[272] = out_r[23:8];
           result_i_ns[272] = out_i[23:8];
        end
        10'd547 : begin
           result_r_ns[784] = out_r[23:8];
           result_i_ns[784] = out_i[23:8];
        end
        10'd548 : begin
           result_r_ns[144] = out_r[23:8];
           result_i_ns[144] = out_i[23:8];
        end
        10'd549 : begin
           result_r_ns[656] = out_r[23:8];
           result_i_ns[656] = out_i[23:8];
        end
        10'd550 : begin
           result_r_ns[400] = out_r[23:8];
           result_i_ns[400] = out_i[23:8];
        end
        10'd551 : begin
           result_r_ns[912] = out_r[23:8];
           result_i_ns[912] = out_i[23:8];
        end
        10'd552 : begin
           result_r_ns[80] = out_r[23:8];
           result_i_ns[80] = out_i[23:8];
        end
        10'd553 : begin
           result_r_ns[592] = out_r[23:8];
           result_i_ns[592] = out_i[23:8];
        end
        10'd554 : begin
           result_r_ns[336] = out_r[23:8];
           result_i_ns[336] = out_i[23:8];
        end
        10'd555 : begin
           result_r_ns[848] = out_r[23:8];
           result_i_ns[848] = out_i[23:8];
        end
        10'd556 : begin
           result_r_ns[208] = out_r[23:8];
           result_i_ns[208] = out_i[23:8];
        end
        10'd557 : begin
           result_r_ns[720] = out_r[23:8];
           result_i_ns[720] = out_i[23:8];
        end
        10'd558 : begin
           result_r_ns[464] = out_r[23:8];
           result_i_ns[464] = out_i[23:8];
        end
        10'd559 : begin
           result_r_ns[976] = out_r[23:8];
           result_i_ns[976] = out_i[23:8];
        end
        10'd560 : begin
           result_r_ns[48] = out_r[23:8];
           result_i_ns[48] = out_i[23:8];
        end
        10'd561 : begin
           result_r_ns[560] = out_r[23:8];
           result_i_ns[560] = out_i[23:8];
        end
        10'd562 : begin
           result_r_ns[304] = out_r[23:8];
           result_i_ns[304] = out_i[23:8];
        end
        10'd563 : begin
           result_r_ns[816] = out_r[23:8];
           result_i_ns[816] = out_i[23:8];
        end
        10'd564 : begin
           result_r_ns[176] = out_r[23:8];
           result_i_ns[176] = out_i[23:8];
        end
        10'd565 : begin
           result_r_ns[688] = out_r[23:8];
           result_i_ns[688] = out_i[23:8];
        end
        10'd566 : begin
           result_r_ns[432] = out_r[23:8];
           result_i_ns[432] = out_i[23:8];
        end
        10'd567 : begin
           result_r_ns[944] = out_r[23:8];
           result_i_ns[944] = out_i[23:8];
        end
        10'd568 : begin
           result_r_ns[112] = out_r[23:8];
           result_i_ns[112] = out_i[23:8];
        end
        10'd569 : begin
           result_r_ns[624] = out_r[23:8];
           result_i_ns[624] = out_i[23:8];
        end
        10'd570 : begin
           result_r_ns[368] = out_r[23:8];
           result_i_ns[368] = out_i[23:8];
        end
        10'd571 : begin
           result_r_ns[880] = out_r[23:8];
           result_i_ns[880] = out_i[23:8];
        end
        10'd572 : begin
           result_r_ns[240] = out_r[23:8];
           result_i_ns[240] = out_i[23:8];
        end
        10'd573 : begin
           result_r_ns[752] = out_r[23:8];
           result_i_ns[752] = out_i[23:8];
        end
        10'd574 : begin
           result_r_ns[496] = out_r[23:8];
           result_i_ns[496] = out_i[23:8];
        end
        10'd575 : begin
           result_r_ns[1008] = out_r[23:8];
           result_i_ns[1008] = out_i[23:8];
        end
        10'd576 : begin
           result_r_ns[8] = out_r[23:8];
           result_i_ns[8] = out_i[23:8];
        end
        10'd577 : begin
           result_r_ns[520] = out_r[23:8];
           result_i_ns[520] = out_i[23:8];
        end
        10'd578 : begin
           result_r_ns[264] = out_r[23:8];
           result_i_ns[264] = out_i[23:8];
        end
        10'd579 : begin
           result_r_ns[776] = out_r[23:8];
           result_i_ns[776] = out_i[23:8];
        end
        10'd580 : begin
           result_r_ns[136] = out_r[23:8];
           result_i_ns[136] = out_i[23:8];
        end
        10'd581 : begin
           result_r_ns[648] = out_r[23:8];
           result_i_ns[648] = out_i[23:8];
        end
        10'd582 : begin
           result_r_ns[392] = out_r[23:8];
           result_i_ns[392] = out_i[23:8];
        end
        10'd583 : begin
           result_r_ns[904] = out_r[23:8];
           result_i_ns[904] = out_i[23:8];
        end
        10'd584 : begin
           result_r_ns[72] = out_r[23:8];
           result_i_ns[72] = out_i[23:8];
        end
        10'd585 : begin
           result_r_ns[584] = out_r[23:8];
           result_i_ns[584] = out_i[23:8];
        end
        10'd586 : begin
           result_r_ns[328] = out_r[23:8];
           result_i_ns[328] = out_i[23:8];
        end
        10'd587 : begin
           result_r_ns[840] = out_r[23:8];
           result_i_ns[840] = out_i[23:8];
        end
        10'd588 : begin
           result_r_ns[200] = out_r[23:8];
           result_i_ns[200] = out_i[23:8];
        end
        10'd589 : begin
           result_r_ns[712] = out_r[23:8];
           result_i_ns[712] = out_i[23:8];
        end
        10'd590 : begin
           result_r_ns[456] = out_r[23:8];
           result_i_ns[456] = out_i[23:8];
        end
        10'd591 : begin
           result_r_ns[968] = out_r[23:8];
           result_i_ns[968] = out_i[23:8];
        end
        10'd592 : begin
           result_r_ns[40] = out_r[23:8];
           result_i_ns[40] = out_i[23:8];
        end
        10'd593 : begin
           result_r_ns[552] = out_r[23:8];
           result_i_ns[552] = out_i[23:8];
        end
        10'd594 : begin
           result_r_ns[296] = out_r[23:8];
           result_i_ns[296] = out_i[23:8];
        end
        10'd595 : begin
           result_r_ns[808] = out_r[23:8];
           result_i_ns[808] = out_i[23:8];
        end
        10'd596 : begin
           result_r_ns[168] = out_r[23:8];
           result_i_ns[168] = out_i[23:8];
        end
        10'd597 : begin
           result_r_ns[680] = out_r[23:8];
           result_i_ns[680] = out_i[23:8];
        end
        10'd598 : begin
           result_r_ns[424] = out_r[23:8];
           result_i_ns[424] = out_i[23:8];
        end
        10'd599 : begin
           result_r_ns[936] = out_r[23:8];
           result_i_ns[936] = out_i[23:8];
        end
        10'd600 : begin
           result_r_ns[104] = out_r[23:8];
           result_i_ns[104] = out_i[23:8];
        end
        10'd601 : begin
           result_r_ns[616] = out_r[23:8];
           result_i_ns[616] = out_i[23:8];
        end
        10'd602 : begin
           result_r_ns[360] = out_r[23:8];
           result_i_ns[360] = out_i[23:8];
        end
        10'd603 : begin
           result_r_ns[872] = out_r[23:8];
           result_i_ns[872] = out_i[23:8];
        end
        10'd604 : begin
           result_r_ns[232] = out_r[23:8];
           result_i_ns[232] = out_i[23:8];
        end
        10'd605 : begin
           result_r_ns[744] = out_r[23:8];
           result_i_ns[744] = out_i[23:8];
        end
        10'd606 : begin
           result_r_ns[488] = out_r[23:8];
           result_i_ns[488] = out_i[23:8];
        end
        10'd607 : begin
           result_r_ns[1000] = out_r[23:8];
           result_i_ns[1000] = out_i[23:8];
        end
        10'd608 : begin
           result_r_ns[24] = out_r[23:8];
           result_i_ns[24] = out_i[23:8];
        end
        10'd609 : begin
           result_r_ns[536] = out_r[23:8];
           result_i_ns[536] = out_i[23:8];
        end
        10'd610 : begin
           result_r_ns[280] = out_r[23:8];
           result_i_ns[280] = out_i[23:8];
        end
        10'd611 : begin
           result_r_ns[792] = out_r[23:8];
           result_i_ns[792] = out_i[23:8];
        end
        10'd612 : begin
           result_r_ns[152] = out_r[23:8];
           result_i_ns[152] = out_i[23:8];
        end
        10'd613 : begin
           result_r_ns[664] = out_r[23:8];
           result_i_ns[664] = out_i[23:8];
        end
        10'd614 : begin
           result_r_ns[408] = out_r[23:8];
           result_i_ns[408] = out_i[23:8];
        end
        10'd615 : begin
           result_r_ns[920] = out_r[23:8];
           result_i_ns[920] = out_i[23:8];
        end
        10'd616 : begin
           result_r_ns[88] = out_r[23:8];
           result_i_ns[88] = out_i[23:8];
        end
        10'd617 : begin
           result_r_ns[600] = out_r[23:8];
           result_i_ns[600] = out_i[23:8];
        end
        10'd618 : begin
           result_r_ns[344] = out_r[23:8];
           result_i_ns[344] = out_i[23:8];
        end
        10'd619 : begin
           result_r_ns[856] = out_r[23:8];
           result_i_ns[856] = out_i[23:8];
        end
        10'd620 : begin
           result_r_ns[216] = out_r[23:8];
           result_i_ns[216] = out_i[23:8];
        end
        10'd621 : begin
           result_r_ns[728] = out_r[23:8];
           result_i_ns[728] = out_i[23:8];
        end
        10'd622 : begin
           result_r_ns[472] = out_r[23:8];
           result_i_ns[472] = out_i[23:8];
        end
        10'd623 : begin
           result_r_ns[984] = out_r[23:8];
           result_i_ns[984] = out_i[23:8];
        end
        10'd624 : begin
           result_r_ns[56] = out_r[23:8];
           result_i_ns[56] = out_i[23:8];
        end
        10'd625 : begin
           result_r_ns[568] = out_r[23:8];
           result_i_ns[568] = out_i[23:8];
        end
        10'd626 : begin
           result_r_ns[312] = out_r[23:8];
           result_i_ns[312] = out_i[23:8];
        end
        10'd627 : begin
           result_r_ns[824] = out_r[23:8];
           result_i_ns[824] = out_i[23:8];
        end
        10'd628 : begin
           result_r_ns[184] = out_r[23:8];
           result_i_ns[184] = out_i[23:8];
        end
        10'd629 : begin
           result_r_ns[696] = out_r[23:8];
           result_i_ns[696] = out_i[23:8];
        end
        10'd630 : begin
           result_r_ns[440] = out_r[23:8];
           result_i_ns[440] = out_i[23:8];
        end
        10'd631 : begin
           result_r_ns[952] = out_r[23:8];
           result_i_ns[952] = out_i[23:8];
        end
        10'd632 : begin
           result_r_ns[120] = out_r[23:8];
           result_i_ns[120] = out_i[23:8];
        end
        10'd633 : begin
           result_r_ns[632] = out_r[23:8];
           result_i_ns[632] = out_i[23:8];
        end
        10'd634 : begin
           result_r_ns[376] = out_r[23:8];
           result_i_ns[376] = out_i[23:8];
        end
        10'd635 : begin
           result_r_ns[888] = out_r[23:8];
           result_i_ns[888] = out_i[23:8];
        end
        10'd636 : begin
           result_r_ns[248] = out_r[23:8];
           result_i_ns[248] = out_i[23:8];
        end
        10'd637 : begin
           result_r_ns[760] = out_r[23:8];
           result_i_ns[760] = out_i[23:8];
        end
        10'd638 : begin
           result_r_ns[504] = out_r[23:8];
           result_i_ns[504] = out_i[23:8];
        end
        10'd639 : begin
           result_r_ns[1016] = out_r[23:8];
           result_i_ns[1016] = out_i[23:8];
        end
        10'd640 : begin
           result_r_ns[4] = out_r[23:8];
           result_i_ns[4] = out_i[23:8];
        end
        10'd641 : begin
           result_r_ns[516] = out_r[23:8];
           result_i_ns[516] = out_i[23:8];
        end
        10'd642 : begin
           result_r_ns[260] = out_r[23:8];
           result_i_ns[260] = out_i[23:8];
        end
        10'd643 : begin
           result_r_ns[772] = out_r[23:8];
           result_i_ns[772] = out_i[23:8];
        end
        10'd644 : begin
           result_r_ns[132] = out_r[23:8];
           result_i_ns[132] = out_i[23:8];
        end
        10'd645 : begin
           result_r_ns[644] = out_r[23:8];
           result_i_ns[644] = out_i[23:8];
        end
        10'd646 : begin
           result_r_ns[388] = out_r[23:8];
           result_i_ns[388] = out_i[23:8];
        end
        10'd647 : begin
           result_r_ns[900] = out_r[23:8];
           result_i_ns[900] = out_i[23:8];
        end
        10'd648 : begin
           result_r_ns[68] = out_r[23:8];
           result_i_ns[68] = out_i[23:8];
        end
        10'd649 : begin
           result_r_ns[580] = out_r[23:8];
           result_i_ns[580] = out_i[23:8];
        end
        10'd650 : begin
           result_r_ns[324] = out_r[23:8];
           result_i_ns[324] = out_i[23:8];
        end
        10'd651 : begin
           result_r_ns[836] = out_r[23:8];
           result_i_ns[836] = out_i[23:8];
        end
        10'd652 : begin
           result_r_ns[196] = out_r[23:8];
           result_i_ns[196] = out_i[23:8];
        end
        10'd653 : begin
           result_r_ns[708] = out_r[23:8];
           result_i_ns[708] = out_i[23:8];
        end
        10'd654 : begin
           result_r_ns[452] = out_r[23:8];
           result_i_ns[452] = out_i[23:8];
        end
        10'd655 : begin
           result_r_ns[964] = out_r[23:8];
           result_i_ns[964] = out_i[23:8];
        end
        10'd656 : begin
           result_r_ns[36] = out_r[23:8];
           result_i_ns[36] = out_i[23:8];
        end
        10'd657 : begin
           result_r_ns[548] = out_r[23:8];
           result_i_ns[548] = out_i[23:8];
        end
        10'd658 : begin
           result_r_ns[292] = out_r[23:8];
           result_i_ns[292] = out_i[23:8];
        end
        10'd659 : begin
           result_r_ns[804] = out_r[23:8];
           result_i_ns[804] = out_i[23:8];
        end
        10'd660 : begin
           result_r_ns[164] = out_r[23:8];
           result_i_ns[164] = out_i[23:8];
        end
        10'd661 : begin
           result_r_ns[676] = out_r[23:8];
           result_i_ns[676] = out_i[23:8];
        end
        10'd662 : begin
           result_r_ns[420] = out_r[23:8];
           result_i_ns[420] = out_i[23:8];
        end
        10'd663 : begin
           result_r_ns[932] = out_r[23:8];
           result_i_ns[932] = out_i[23:8];
        end
        10'd664 : begin
           result_r_ns[100] = out_r[23:8];
           result_i_ns[100] = out_i[23:8];
        end
        10'd665 : begin
           result_r_ns[612] = out_r[23:8];
           result_i_ns[612] = out_i[23:8];
        end
        10'd666 : begin
           result_r_ns[356] = out_r[23:8];
           result_i_ns[356] = out_i[23:8];
        end
        10'd667 : begin
           result_r_ns[868] = out_r[23:8];
           result_i_ns[868] = out_i[23:8];
        end
        10'd668 : begin
           result_r_ns[228] = out_r[23:8];
           result_i_ns[228] = out_i[23:8];
        end
        10'd669 : begin
           result_r_ns[740] = out_r[23:8];
           result_i_ns[740] = out_i[23:8];
        end
        10'd670 : begin
           result_r_ns[484] = out_r[23:8];
           result_i_ns[484] = out_i[23:8];
        end
        10'd671 : begin
           result_r_ns[996] = out_r[23:8];
           result_i_ns[996] = out_i[23:8];
        end
        10'd672 : begin
           result_r_ns[20] = out_r[23:8];
           result_i_ns[20] = out_i[23:8];
        end
        10'd673 : begin
           result_r_ns[532] = out_r[23:8];
           result_i_ns[532] = out_i[23:8];
        end
        10'd674 : begin
           result_r_ns[276] = out_r[23:8];
           result_i_ns[276] = out_i[23:8];
        end
        10'd675 : begin
           result_r_ns[788] = out_r[23:8];
           result_i_ns[788] = out_i[23:8];
        end
        10'd676 : begin
           result_r_ns[148] = out_r[23:8];
           result_i_ns[148] = out_i[23:8];
        end
        10'd677 : begin
           result_r_ns[660] = out_r[23:8];
           result_i_ns[660] = out_i[23:8];
        end
        10'd678 : begin
           result_r_ns[404] = out_r[23:8];
           result_i_ns[404] = out_i[23:8];
        end
        10'd679 : begin
           result_r_ns[916] = out_r[23:8];
           result_i_ns[916] = out_i[23:8];
        end
        10'd680 : begin
           result_r_ns[84] = out_r[23:8];
           result_i_ns[84] = out_i[23:8];
        end
        10'd681 : begin
           result_r_ns[596] = out_r[23:8];
           result_i_ns[596] = out_i[23:8];
        end
        10'd682 : begin
           result_r_ns[340] = out_r[23:8];
           result_i_ns[340] = out_i[23:8];
        end
        10'd683 : begin
           result_r_ns[852] = out_r[23:8];
           result_i_ns[852] = out_i[23:8];
        end
        10'd684 : begin
           result_r_ns[212] = out_r[23:8];
           result_i_ns[212] = out_i[23:8];
        end
        10'd685 : begin
           result_r_ns[724] = out_r[23:8];
           result_i_ns[724] = out_i[23:8];
        end
        10'd686 : begin
           result_r_ns[468] = out_r[23:8];
           result_i_ns[468] = out_i[23:8];
        end
        10'd687 : begin
           result_r_ns[980] = out_r[23:8];
           result_i_ns[980] = out_i[23:8];
        end
        10'd688 : begin
           result_r_ns[52] = out_r[23:8];
           result_i_ns[52] = out_i[23:8];
        end
        10'd689 : begin
           result_r_ns[564] = out_r[23:8];
           result_i_ns[564] = out_i[23:8];
        end
        10'd690 : begin
           result_r_ns[308] = out_r[23:8];
           result_i_ns[308] = out_i[23:8];
        end
        10'd691 : begin
           result_r_ns[820] = out_r[23:8];
           result_i_ns[820] = out_i[23:8];
        end
        10'd692 : begin
           result_r_ns[180] = out_r[23:8];
           result_i_ns[180] = out_i[23:8];
        end
        10'd693 : begin
           result_r_ns[692] = out_r[23:8];
           result_i_ns[692] = out_i[23:8];
        end
        10'd694 : begin
           result_r_ns[436] = out_r[23:8];
           result_i_ns[436] = out_i[23:8];
        end
        10'd695 : begin
           result_r_ns[948] = out_r[23:8];
           result_i_ns[948] = out_i[23:8];
        end
        10'd696 : begin
           result_r_ns[116] = out_r[23:8];
           result_i_ns[116] = out_i[23:8];
        end
        10'd697 : begin
           result_r_ns[628] = out_r[23:8];
           result_i_ns[628] = out_i[23:8];
        end
        10'd698 : begin
           result_r_ns[372] = out_r[23:8];
           result_i_ns[372] = out_i[23:8];
        end
        10'd699 : begin
           result_r_ns[884] = out_r[23:8];
           result_i_ns[884] = out_i[23:8];
        end
        10'd700 : begin
           result_r_ns[244] = out_r[23:8];
           result_i_ns[244] = out_i[23:8];
        end
        10'd701 : begin
           result_r_ns[756] = out_r[23:8];
           result_i_ns[756] = out_i[23:8];
        end
        10'd702 : begin
           result_r_ns[500] = out_r[23:8];
           result_i_ns[500] = out_i[23:8];
        end
        10'd703 : begin
           result_r_ns[1012] = out_r[23:8];
           result_i_ns[1012] = out_i[23:8];
        end
        10'd704 : begin
           result_r_ns[12] = out_r[23:8];
           result_i_ns[12] = out_i[23:8];
        end
        10'd705 : begin
           result_r_ns[524] = out_r[23:8];
           result_i_ns[524] = out_i[23:8];
        end
        10'd706 : begin
           result_r_ns[268] = out_r[23:8];
           result_i_ns[268] = out_i[23:8];
        end
        10'd707 : begin
           result_r_ns[780] = out_r[23:8];
           result_i_ns[780] = out_i[23:8];
        end
        10'd708 : begin
           result_r_ns[140] = out_r[23:8];
           result_i_ns[140] = out_i[23:8];
        end
        10'd709 : begin
           result_r_ns[652] = out_r[23:8];
           result_i_ns[652] = out_i[23:8];
        end
        10'd710 : begin
           result_r_ns[396] = out_r[23:8];
           result_i_ns[396] = out_i[23:8];
        end
        10'd711 : begin
           result_r_ns[908] = out_r[23:8];
           result_i_ns[908] = out_i[23:8];
        end
        10'd712 : begin
           result_r_ns[76] = out_r[23:8];
           result_i_ns[76] = out_i[23:8];
        end
        10'd713 : begin
           result_r_ns[588] = out_r[23:8];
           result_i_ns[588] = out_i[23:8];
        end
        10'd714 : begin
           result_r_ns[332] = out_r[23:8];
           result_i_ns[332] = out_i[23:8];
        end
        10'd715 : begin
           result_r_ns[844] = out_r[23:8];
           result_i_ns[844] = out_i[23:8];
        end
        10'd716 : begin
           result_r_ns[204] = out_r[23:8];
           result_i_ns[204] = out_i[23:8];
        end
        10'd717 : begin
           result_r_ns[716] = out_r[23:8];
           result_i_ns[716] = out_i[23:8];
        end
        10'd718 : begin
           result_r_ns[460] = out_r[23:8];
           result_i_ns[460] = out_i[23:8];
        end
        10'd719 : begin
           result_r_ns[972] = out_r[23:8];
           result_i_ns[972] = out_i[23:8];
        end
        10'd720 : begin
           result_r_ns[44] = out_r[23:8];
           result_i_ns[44] = out_i[23:8];
        end
        10'd721 : begin
           result_r_ns[556] = out_r[23:8];
           result_i_ns[556] = out_i[23:8];
        end
        10'd722 : begin
           result_r_ns[300] = out_r[23:8];
           result_i_ns[300] = out_i[23:8];
        end
        10'd723 : begin
           result_r_ns[812] = out_r[23:8];
           result_i_ns[812] = out_i[23:8];
        end
        10'd724 : begin
           result_r_ns[172] = out_r[23:8];
           result_i_ns[172] = out_i[23:8];
        end
        10'd725 : begin
           result_r_ns[684] = out_r[23:8];
           result_i_ns[684] = out_i[23:8];
        end
        10'd726 : begin
           result_r_ns[428] = out_r[23:8];
           result_i_ns[428] = out_i[23:8];
        end
        10'd727 : begin
           result_r_ns[940] = out_r[23:8];
           result_i_ns[940] = out_i[23:8];
        end
        10'd728 : begin
           result_r_ns[108] = out_r[23:8];
           result_i_ns[108] = out_i[23:8];
        end
        10'd729 : begin
           result_r_ns[620] = out_r[23:8];
           result_i_ns[620] = out_i[23:8];
        end
        10'd730 : begin
           result_r_ns[364] = out_r[23:8];
           result_i_ns[364] = out_i[23:8];
        end
        10'd731 : begin
           result_r_ns[876] = out_r[23:8];
           result_i_ns[876] = out_i[23:8];
        end
        10'd732 : begin
           result_r_ns[236] = out_r[23:8];
           result_i_ns[236] = out_i[23:8];
        end
        10'd733 : begin
           result_r_ns[748] = out_r[23:8];
           result_i_ns[748] = out_i[23:8];
        end
        10'd734 : begin
           result_r_ns[492] = out_r[23:8];
           result_i_ns[492] = out_i[23:8];
        end
        10'd735 : begin
           result_r_ns[1004] = out_r[23:8];
           result_i_ns[1004] = out_i[23:8];
        end
        10'd736 : begin
           result_r_ns[28] = out_r[23:8];
           result_i_ns[28] = out_i[23:8];
        end
        10'd737 : begin
           result_r_ns[540] = out_r[23:8];
           result_i_ns[540] = out_i[23:8];
        end
        10'd738 : begin
           result_r_ns[284] = out_r[23:8];
           result_i_ns[284] = out_i[23:8];
        end
        10'd739 : begin
           result_r_ns[796] = out_r[23:8];
           result_i_ns[796] = out_i[23:8];
        end
        10'd740 : begin
           result_r_ns[156] = out_r[23:8];
           result_i_ns[156] = out_i[23:8];
        end
        10'd741 : begin
           result_r_ns[668] = out_r[23:8];
           result_i_ns[668] = out_i[23:8];
        end
        10'd742 : begin
           result_r_ns[412] = out_r[23:8];
           result_i_ns[412] = out_i[23:8];
        end
        10'd743 : begin
           result_r_ns[924] = out_r[23:8];
           result_i_ns[924] = out_i[23:8];
        end
        10'd744 : begin
           result_r_ns[92] = out_r[23:8];
           result_i_ns[92] = out_i[23:8];
        end
        10'd745 : begin
           result_r_ns[604] = out_r[23:8];
           result_i_ns[604] = out_i[23:8];
        end
        10'd746 : begin
           result_r_ns[348] = out_r[23:8];
           result_i_ns[348] = out_i[23:8];
        end
        10'd747 : begin
           result_r_ns[860] = out_r[23:8];
           result_i_ns[860] = out_i[23:8];
        end
        10'd748 : begin
           result_r_ns[220] = out_r[23:8];
           result_i_ns[220] = out_i[23:8];
        end
        10'd749 : begin
           result_r_ns[732] = out_r[23:8];
           result_i_ns[732] = out_i[23:8];
        end
        10'd750 : begin
           result_r_ns[476] = out_r[23:8];
           result_i_ns[476] = out_i[23:8];
        end
        10'd751 : begin
           result_r_ns[988] = out_r[23:8];
           result_i_ns[988] = out_i[23:8];
        end
        10'd752 : begin
           result_r_ns[60] = out_r[23:8];
           result_i_ns[60] = out_i[23:8];
        end
        10'd753 : begin
           result_r_ns[572] = out_r[23:8];
           result_i_ns[572] = out_i[23:8];
        end
        10'd754 : begin
           result_r_ns[316] = out_r[23:8];
           result_i_ns[316] = out_i[23:8];
        end
        10'd755 : begin
           result_r_ns[828] = out_r[23:8];
           result_i_ns[828] = out_i[23:8];
        end
        10'd756 : begin
           result_r_ns[188] = out_r[23:8];
           result_i_ns[188] = out_i[23:8];
        end
        10'd757 : begin
           result_r_ns[700] = out_r[23:8];
           result_i_ns[700] = out_i[23:8];
        end
        10'd758 : begin
           result_r_ns[444] = out_r[23:8];
           result_i_ns[444] = out_i[23:8];
        end
        10'd759 : begin
           result_r_ns[956] = out_r[23:8];
           result_i_ns[956] = out_i[23:8];
        end
        10'd760 : begin
           result_r_ns[124] = out_r[23:8];
           result_i_ns[124] = out_i[23:8];
        end
        10'd761 : begin
           result_r_ns[636] = out_r[23:8];
           result_i_ns[636] = out_i[23:8];
        end
        10'd762 : begin
           result_r_ns[380] = out_r[23:8];
           result_i_ns[380] = out_i[23:8];
        end
        10'd763 : begin
           result_r_ns[892] = out_r[23:8];
           result_i_ns[892] = out_i[23:8];
        end
        10'd764 : begin
           result_r_ns[252] = out_r[23:8];
           result_i_ns[252] = out_i[23:8];
        end
        10'd765 : begin
           result_r_ns[764] = out_r[23:8];
           result_i_ns[764] = out_i[23:8];
        end
        10'd766 : begin
           result_r_ns[508] = out_r[23:8];
           result_i_ns[508] = out_i[23:8];
        end
        10'd767 : begin
           result_r_ns[1020] = out_r[23:8];
           result_i_ns[1020] = out_i[23:8];
        end
        10'd768 : begin
           result_r_ns[2] = out_r[23:8];
           result_i_ns[2] = out_i[23:8];
        end
        10'd769 : begin
           result_r_ns[514] = out_r[23:8];
           result_i_ns[514] = out_i[23:8];
        end
        10'd770 : begin
           result_r_ns[258] = out_r[23:8];
           result_i_ns[258] = out_i[23:8];
        end
        10'd771 : begin
           result_r_ns[770] = out_r[23:8];
           result_i_ns[770] = out_i[23:8];
        end
        10'd772 : begin
           result_r_ns[130] = out_r[23:8];
           result_i_ns[130] = out_i[23:8];
        end
        10'd773 : begin
           result_r_ns[642] = out_r[23:8];
           result_i_ns[642] = out_i[23:8];
        end
        10'd774 : begin
           result_r_ns[386] = out_r[23:8];
           result_i_ns[386] = out_i[23:8];
        end
        10'd775 : begin
           result_r_ns[898] = out_r[23:8];
           result_i_ns[898] = out_i[23:8];
        end
        10'd776 : begin
           result_r_ns[66] = out_r[23:8];
           result_i_ns[66] = out_i[23:8];
        end
        10'd777 : begin
           result_r_ns[578] = out_r[23:8];
           result_i_ns[578] = out_i[23:8];
        end
        10'd778 : begin
           result_r_ns[322] = out_r[23:8];
           result_i_ns[322] = out_i[23:8];
        end
        10'd779 : begin
           result_r_ns[834] = out_r[23:8];
           result_i_ns[834] = out_i[23:8];
        end
        10'd780 : begin
           result_r_ns[194] = out_r[23:8];
           result_i_ns[194] = out_i[23:8];
        end
        10'd781 : begin
           result_r_ns[706] = out_r[23:8];
           result_i_ns[706] = out_i[23:8];
        end
        10'd782 : begin
           result_r_ns[450] = out_r[23:8];
           result_i_ns[450] = out_i[23:8];
        end
        10'd783 : begin
           result_r_ns[962] = out_r[23:8];
           result_i_ns[962] = out_i[23:8];
        end
        10'd784 : begin
           result_r_ns[34] = out_r[23:8];
           result_i_ns[34] = out_i[23:8];
        end
        10'd785 : begin
           result_r_ns[546] = out_r[23:8];
           result_i_ns[546] = out_i[23:8];
        end
        10'd786 : begin
           result_r_ns[290] = out_r[23:8];
           result_i_ns[290] = out_i[23:8];
        end
        10'd787 : begin
           result_r_ns[802] = out_r[23:8];
           result_i_ns[802] = out_i[23:8];
        end
        10'd788 : begin
           result_r_ns[162] = out_r[23:8];
           result_i_ns[162] = out_i[23:8];
        end
        10'd789 : begin
           result_r_ns[674] = out_r[23:8];
           result_i_ns[674] = out_i[23:8];
        end
        10'd790 : begin
           result_r_ns[418] = out_r[23:8];
           result_i_ns[418] = out_i[23:8];
        end
        10'd791 : begin
           result_r_ns[930] = out_r[23:8];
           result_i_ns[930] = out_i[23:8];
        end
        10'd792 : begin
           result_r_ns[98] = out_r[23:8];
           result_i_ns[98] = out_i[23:8];
        end
        10'd793 : begin
           result_r_ns[610] = out_r[23:8];
           result_i_ns[610] = out_i[23:8];
        end
        10'd794 : begin
           result_r_ns[354] = out_r[23:8];
           result_i_ns[354] = out_i[23:8];
        end
        10'd795 : begin
           result_r_ns[866] = out_r[23:8];
           result_i_ns[866] = out_i[23:8];
        end
        10'd796 : begin
           result_r_ns[226] = out_r[23:8];
           result_i_ns[226] = out_i[23:8];
        end
        10'd797 : begin
           result_r_ns[738] = out_r[23:8];
           result_i_ns[738] = out_i[23:8];
        end
        10'd798 : begin
           result_r_ns[482] = out_r[23:8];
           result_i_ns[482] = out_i[23:8];
        end
        10'd799 : begin
           result_r_ns[994] = out_r[23:8];
           result_i_ns[994] = out_i[23:8];
        end
        10'd800 : begin
           result_r_ns[18] = out_r[23:8];
           result_i_ns[18] = out_i[23:8];
        end
        10'd801 : begin
           result_r_ns[530] = out_r[23:8];
           result_i_ns[530] = out_i[23:8];
        end
        10'd802 : begin
           result_r_ns[274] = out_r[23:8];
           result_i_ns[274] = out_i[23:8];
        end
        10'd803 : begin
           result_r_ns[786] = out_r[23:8];
           result_i_ns[786] = out_i[23:8];
        end
        10'd804 : begin
           result_r_ns[146] = out_r[23:8];
           result_i_ns[146] = out_i[23:8];
        end
        10'd805 : begin
           result_r_ns[658] = out_r[23:8];
           result_i_ns[658] = out_i[23:8];
        end
        10'd806 : begin
           result_r_ns[402] = out_r[23:8];
           result_i_ns[402] = out_i[23:8];
        end
        10'd807 : begin
           result_r_ns[914] = out_r[23:8];
           result_i_ns[914] = out_i[23:8];
        end
        10'd808 : begin
           result_r_ns[82] = out_r[23:8];
           result_i_ns[82] = out_i[23:8];
        end
        10'd809 : begin
           result_r_ns[594] = out_r[23:8];
           result_i_ns[594] = out_i[23:8];
        end
        10'd810 : begin
           result_r_ns[338] = out_r[23:8];
           result_i_ns[338] = out_i[23:8];
        end
        10'd811 : begin
           result_r_ns[850] = out_r[23:8];
           result_i_ns[850] = out_i[23:8];
        end
        10'd812 : begin
           result_r_ns[210] = out_r[23:8];
           result_i_ns[210] = out_i[23:8];
        end
        10'd813 : begin
           result_r_ns[722] = out_r[23:8];
           result_i_ns[722] = out_i[23:8];
        end
        10'd814 : begin
           result_r_ns[466] = out_r[23:8];
           result_i_ns[466] = out_i[23:8];
        end
        10'd815 : begin
           result_r_ns[978] = out_r[23:8];
           result_i_ns[978] = out_i[23:8];
        end
        10'd816 : begin
           result_r_ns[50] = out_r[23:8];
           result_i_ns[50] = out_i[23:8];
        end
        10'd817 : begin
           result_r_ns[562] = out_r[23:8];
           result_i_ns[562] = out_i[23:8];
        end
        10'd818 : begin
           result_r_ns[306] = out_r[23:8];
           result_i_ns[306] = out_i[23:8];
        end
        10'd819 : begin
           result_r_ns[818] = out_r[23:8];
           result_i_ns[818] = out_i[23:8];
        end
        10'd820 : begin
           result_r_ns[178] = out_r[23:8];
           result_i_ns[178] = out_i[23:8];
        end
        10'd821 : begin
           result_r_ns[690] = out_r[23:8];
           result_i_ns[690] = out_i[23:8];
        end
        10'd822 : begin
           result_r_ns[434] = out_r[23:8];
           result_i_ns[434] = out_i[23:8];
        end
        10'd823 : begin
           result_r_ns[946] = out_r[23:8];
           result_i_ns[946] = out_i[23:8];
        end
        10'd824 : begin
           result_r_ns[114] = out_r[23:8];
           result_i_ns[114] = out_i[23:8];
        end
        10'd825 : begin
           result_r_ns[626] = out_r[23:8];
           result_i_ns[626] = out_i[23:8];
        end
        10'd826 : begin
           result_r_ns[370] = out_r[23:8];
           result_i_ns[370] = out_i[23:8];
        end
        10'd827 : begin
           result_r_ns[882] = out_r[23:8];
           result_i_ns[882] = out_i[23:8];
        end
        10'd828 : begin
           result_r_ns[242] = out_r[23:8];
           result_i_ns[242] = out_i[23:8];
        end
        10'd829 : begin
           result_r_ns[754] = out_r[23:8];
           result_i_ns[754] = out_i[23:8];
        end
        10'd830 : begin
           result_r_ns[498] = out_r[23:8];
           result_i_ns[498] = out_i[23:8];
        end
        10'd831 : begin
           result_r_ns[1010] = out_r[23:8];
           result_i_ns[1010] = out_i[23:8];
        end
        10'd832 : begin
           result_r_ns[10] = out_r[23:8];
           result_i_ns[10] = out_i[23:8];
        end
        10'd833 : begin
           result_r_ns[522] = out_r[23:8];
           result_i_ns[522] = out_i[23:8];
        end
        10'd834 : begin
           result_r_ns[266] = out_r[23:8];
           result_i_ns[266] = out_i[23:8];
        end
        10'd835 : begin
           result_r_ns[778] = out_r[23:8];
           result_i_ns[778] = out_i[23:8];
        end
        10'd836 : begin
           result_r_ns[138] = out_r[23:8];
           result_i_ns[138] = out_i[23:8];
        end
        10'd837 : begin
           result_r_ns[650] = out_r[23:8];
           result_i_ns[650] = out_i[23:8];
        end
        10'd838 : begin
           result_r_ns[394] = out_r[23:8];
           result_i_ns[394] = out_i[23:8];
        end
        10'd839 : begin
           result_r_ns[906] = out_r[23:8];
           result_i_ns[906] = out_i[23:8];
        end
        10'd840 : begin
           result_r_ns[74] = out_r[23:8];
           result_i_ns[74] = out_i[23:8];
        end
        10'd841 : begin
           result_r_ns[586] = out_r[23:8];
           result_i_ns[586] = out_i[23:8];
        end
        10'd842 : begin
           result_r_ns[330] = out_r[23:8];
           result_i_ns[330] = out_i[23:8];
        end
        10'd843 : begin
           result_r_ns[842] = out_r[23:8];
           result_i_ns[842] = out_i[23:8];
        end
        10'd844 : begin
           result_r_ns[202] = out_r[23:8];
           result_i_ns[202] = out_i[23:8];
        end
        10'd845 : begin
           result_r_ns[714] = out_r[23:8];
           result_i_ns[714] = out_i[23:8];
        end
        10'd846 : begin
           result_r_ns[458] = out_r[23:8];
           result_i_ns[458] = out_i[23:8];
        end
        10'd847 : begin
           result_r_ns[970] = out_r[23:8];
           result_i_ns[970] = out_i[23:8];
        end
        10'd848 : begin
           result_r_ns[42] = out_r[23:8];
           result_i_ns[42] = out_i[23:8];
        end
        10'd849 : begin
           result_r_ns[554] = out_r[23:8];
           result_i_ns[554] = out_i[23:8];
        end
        10'd850 : begin
           result_r_ns[298] = out_r[23:8];
           result_i_ns[298] = out_i[23:8];
        end
        10'd851 : begin
           result_r_ns[810] = out_r[23:8];
           result_i_ns[810] = out_i[23:8];
        end
        10'd852 : begin
           result_r_ns[170] = out_r[23:8];
           result_i_ns[170] = out_i[23:8];
        end
        10'd853 : begin
           result_r_ns[682] = out_r[23:8];
           result_i_ns[682] = out_i[23:8];
        end
        10'd854 : begin
           result_r_ns[426] = out_r[23:8];
           result_i_ns[426] = out_i[23:8];
        end
        10'd855 : begin
           result_r_ns[938] = out_r[23:8];
           result_i_ns[938] = out_i[23:8];
        end
        10'd856 : begin
           result_r_ns[106] = out_r[23:8];
           result_i_ns[106] = out_i[23:8];
        end
        10'd857 : begin
           result_r_ns[618] = out_r[23:8];
           result_i_ns[618] = out_i[23:8];
        end
        10'd858 : begin
           result_r_ns[362] = out_r[23:8];
           result_i_ns[362] = out_i[23:8];
        end
        10'd859 : begin
           result_r_ns[874] = out_r[23:8];
           result_i_ns[874] = out_i[23:8];
        end
        10'd860 : begin
           result_r_ns[234] = out_r[23:8];
           result_i_ns[234] = out_i[23:8];
        end
        10'd861 : begin
           result_r_ns[746] = out_r[23:8];
           result_i_ns[746] = out_i[23:8];
        end
        10'd862 : begin
           result_r_ns[490] = out_r[23:8];
           result_i_ns[490] = out_i[23:8];
        end
        10'd863 : begin
           result_r_ns[1002] = out_r[23:8];
           result_i_ns[1002] = out_i[23:8];
        end
        10'd864 : begin
           result_r_ns[26] = out_r[23:8];
           result_i_ns[26] = out_i[23:8];
        end
        10'd865 : begin
           result_r_ns[538] = out_r[23:8];
           result_i_ns[538] = out_i[23:8];
        end
        10'd866 : begin
           result_r_ns[282] = out_r[23:8];
           result_i_ns[282] = out_i[23:8];
        end
        10'd867 : begin
           result_r_ns[794] = out_r[23:8];
           result_i_ns[794] = out_i[23:8];
        end
        10'd868 : begin
           result_r_ns[154] = out_r[23:8];
           result_i_ns[154] = out_i[23:8];
        end
        10'd869 : begin
           result_r_ns[666] = out_r[23:8];
           result_i_ns[666] = out_i[23:8];
        end
        10'd870 : begin
           result_r_ns[410] = out_r[23:8];
           result_i_ns[410] = out_i[23:8];
        end
        10'd871 : begin
           result_r_ns[922] = out_r[23:8];
           result_i_ns[922] = out_i[23:8];
        end
        10'd872 : begin
           result_r_ns[90] = out_r[23:8];
           result_i_ns[90] = out_i[23:8];
        end
        10'd873 : begin
           result_r_ns[602] = out_r[23:8];
           result_i_ns[602] = out_i[23:8];
        end
        10'd874 : begin
           result_r_ns[346] = out_r[23:8];
           result_i_ns[346] = out_i[23:8];
        end
        10'd875 : begin
           result_r_ns[858] = out_r[23:8];
           result_i_ns[858] = out_i[23:8];
        end
        10'd876 : begin
           result_r_ns[218] = out_r[23:8];
           result_i_ns[218] = out_i[23:8];
        end
        10'd877 : begin
           result_r_ns[730] = out_r[23:8];
           result_i_ns[730] = out_i[23:8];
        end
        10'd878 : begin
           result_r_ns[474] = out_r[23:8];
           result_i_ns[474] = out_i[23:8];
        end
        10'd879 : begin
           result_r_ns[986] = out_r[23:8];
           result_i_ns[986] = out_i[23:8];
        end
        10'd880 : begin
           result_r_ns[58] = out_r[23:8];
           result_i_ns[58] = out_i[23:8];
        end
        10'd881 : begin
           result_r_ns[570] = out_r[23:8];
           result_i_ns[570] = out_i[23:8];
        end
        10'd882 : begin
           result_r_ns[314] = out_r[23:8];
           result_i_ns[314] = out_i[23:8];
        end
        10'd883 : begin
           result_r_ns[826] = out_r[23:8];
           result_i_ns[826] = out_i[23:8];
        end
        10'd884 : begin
           result_r_ns[186] = out_r[23:8];
           result_i_ns[186] = out_i[23:8];
        end
        10'd885 : begin
           result_r_ns[698] = out_r[23:8];
           result_i_ns[698] = out_i[23:8];
        end
        10'd886 : begin
           result_r_ns[442] = out_r[23:8];
           result_i_ns[442] = out_i[23:8];
        end
        10'd887 : begin
           result_r_ns[954] = out_r[23:8];
           result_i_ns[954] = out_i[23:8];
        end
        10'd888 : begin
           result_r_ns[122] = out_r[23:8];
           result_i_ns[122] = out_i[23:8];
        end
        10'd889 : begin
           result_r_ns[634] = out_r[23:8];
           result_i_ns[634] = out_i[23:8];
        end
        10'd890 : begin
           result_r_ns[378] = out_r[23:8];
           result_i_ns[378] = out_i[23:8];
        end
        10'd891 : begin
           result_r_ns[890] = out_r[23:8];
           result_i_ns[890] = out_i[23:8];
        end
        10'd892 : begin
           result_r_ns[250] = out_r[23:8];
           result_i_ns[250] = out_i[23:8];
        end
        10'd893 : begin
           result_r_ns[762] = out_r[23:8];
           result_i_ns[762] = out_i[23:8];
        end
        10'd894 : begin
           result_r_ns[506] = out_r[23:8];
           result_i_ns[506] = out_i[23:8];
        end
        10'd895 : begin
           result_r_ns[1018] = out_r[23:8];
           result_i_ns[1018] = out_i[23:8];
        end
        10'd896 : begin
           result_r_ns[6] = out_r[23:8];
           result_i_ns[6] = out_i[23:8];
        end
        10'd897 : begin
           result_r_ns[518] = out_r[23:8];
           result_i_ns[518] = out_i[23:8];
        end
        10'd898 : begin
           result_r_ns[262] = out_r[23:8];
           result_i_ns[262] = out_i[23:8];
        end
        10'd899 : begin
           result_r_ns[774] = out_r[23:8];
           result_i_ns[774] = out_i[23:8];
        end
        10'd900 : begin
           result_r_ns[134] = out_r[23:8];
           result_i_ns[134] = out_i[23:8];
        end
        10'd901 : begin
           result_r_ns[646] = out_r[23:8];
           result_i_ns[646] = out_i[23:8];
        end
        10'd902 : begin
           result_r_ns[390] = out_r[23:8];
           result_i_ns[390] = out_i[23:8];
        end
        10'd903 : begin
           result_r_ns[902] = out_r[23:8];
           result_i_ns[902] = out_i[23:8];
        end
        10'd904 : begin
           result_r_ns[70] = out_r[23:8];
           result_i_ns[70] = out_i[23:8];
        end
        10'd905 : begin
           result_r_ns[582] = out_r[23:8];
           result_i_ns[582] = out_i[23:8];
        end
        10'd906 : begin
           result_r_ns[326] = out_r[23:8];
           result_i_ns[326] = out_i[23:8];
        end
        10'd907 : begin
           result_r_ns[838] = out_r[23:8];
           result_i_ns[838] = out_i[23:8];
        end
        10'd908 : begin
           result_r_ns[198] = out_r[23:8];
           result_i_ns[198] = out_i[23:8];
        end
        10'd909 : begin
           result_r_ns[710] = out_r[23:8];
           result_i_ns[710] = out_i[23:8];
        end
        10'd910 : begin
           result_r_ns[454] = out_r[23:8];
           result_i_ns[454] = out_i[23:8];
        end
        10'd911 : begin
           result_r_ns[966] = out_r[23:8];
           result_i_ns[966] = out_i[23:8];
        end
        10'd912 : begin
           result_r_ns[38] = out_r[23:8];
           result_i_ns[38] = out_i[23:8];
        end
        10'd913 : begin
           result_r_ns[550] = out_r[23:8];
           result_i_ns[550] = out_i[23:8];
        end
        10'd914 : begin
           result_r_ns[294] = out_r[23:8];
           result_i_ns[294] = out_i[23:8];
        end
        10'd915 : begin
           result_r_ns[806] = out_r[23:8];
           result_i_ns[806] = out_i[23:8];
        end
        10'd916 : begin
           result_r_ns[166] = out_r[23:8];
           result_i_ns[166] = out_i[23:8];
        end
        10'd917 : begin
           result_r_ns[678] = out_r[23:8];
           result_i_ns[678] = out_i[23:8];
        end
        10'd918 : begin
           result_r_ns[422] = out_r[23:8];
           result_i_ns[422] = out_i[23:8];
        end
        10'd919 : begin
           result_r_ns[934] = out_r[23:8];
           result_i_ns[934] = out_i[23:8];
        end
        10'd920 : begin
           result_r_ns[102] = out_r[23:8];
           result_i_ns[102] = out_i[23:8];
        end
        10'd921 : begin
           result_r_ns[614] = out_r[23:8];
           result_i_ns[614] = out_i[23:8];
        end
        10'd922 : begin
           result_r_ns[358] = out_r[23:8];
           result_i_ns[358] = out_i[23:8];
        end
        10'd923 : begin
           result_r_ns[870] = out_r[23:8];
           result_i_ns[870] = out_i[23:8];
        end
        10'd924 : begin
           result_r_ns[230] = out_r[23:8];
           result_i_ns[230] = out_i[23:8];
        end
        10'd925 : begin
           result_r_ns[742] = out_r[23:8];
           result_i_ns[742] = out_i[23:8];
        end
        10'd926 : begin
           result_r_ns[486] = out_r[23:8];
           result_i_ns[486] = out_i[23:8];
        end
        10'd927 : begin
           result_r_ns[998] = out_r[23:8];
           result_i_ns[998] = out_i[23:8];
        end
        10'd928 : begin
           result_r_ns[22] = out_r[23:8];
           result_i_ns[22] = out_i[23:8];
        end
        10'd929 : begin
           result_r_ns[534] = out_r[23:8];
           result_i_ns[534] = out_i[23:8];
        end
        10'd930 : begin
           result_r_ns[278] = out_r[23:8];
           result_i_ns[278] = out_i[23:8];
        end
        10'd931 : begin
           result_r_ns[790] = out_r[23:8];
           result_i_ns[790] = out_i[23:8];
        end
        10'd932 : begin
           result_r_ns[150] = out_r[23:8];
           result_i_ns[150] = out_i[23:8];
        end
        10'd933 : begin
           result_r_ns[662] = out_r[23:8];
           result_i_ns[662] = out_i[23:8];
        end
        10'd934 : begin
           result_r_ns[406] = out_r[23:8];
           result_i_ns[406] = out_i[23:8];
        end
        10'd935 : begin
           result_r_ns[918] = out_r[23:8];
           result_i_ns[918] = out_i[23:8];
        end
        10'd936 : begin
           result_r_ns[86] = out_r[23:8];
           result_i_ns[86] = out_i[23:8];
        end
        10'd937 : begin
           result_r_ns[598] = out_r[23:8];
           result_i_ns[598] = out_i[23:8];
        end
        10'd938 : begin
           result_r_ns[342] = out_r[23:8];
           result_i_ns[342] = out_i[23:8];
        end
        10'd939 : begin
           result_r_ns[854] = out_r[23:8];
           result_i_ns[854] = out_i[23:8];
        end
        10'd940 : begin
           result_r_ns[214] = out_r[23:8];
           result_i_ns[214] = out_i[23:8];
        end
        10'd941 : begin
           result_r_ns[726] = out_r[23:8];
           result_i_ns[726] = out_i[23:8];
        end
        10'd942 : begin
           result_r_ns[470] = out_r[23:8];
           result_i_ns[470] = out_i[23:8];
        end
        10'd943 : begin
           result_r_ns[982] = out_r[23:8];
           result_i_ns[982] = out_i[23:8];
        end
        10'd944 : begin
           result_r_ns[54] = out_r[23:8];
           result_i_ns[54] = out_i[23:8];
        end
        10'd945 : begin
           result_r_ns[566] = out_r[23:8];
           result_i_ns[566] = out_i[23:8];
        end
        10'd946 : begin
           result_r_ns[310] = out_r[23:8];
           result_i_ns[310] = out_i[23:8];
        end
        10'd947 : begin
           result_r_ns[822] = out_r[23:8];
           result_i_ns[822] = out_i[23:8];
        end
        10'd948 : begin
           result_r_ns[182] = out_r[23:8];
           result_i_ns[182] = out_i[23:8];
        end
        10'd949 : begin
           result_r_ns[694] = out_r[23:8];
           result_i_ns[694] = out_i[23:8];
        end
        10'd950 : begin
           result_r_ns[438] = out_r[23:8];
           result_i_ns[438] = out_i[23:8];
        end
        10'd951 : begin
           result_r_ns[950] = out_r[23:8];
           result_i_ns[950] = out_i[23:8];
        end
        10'd952 : begin
           result_r_ns[118] = out_r[23:8];
           result_i_ns[118] = out_i[23:8];
        end
        10'd953 : begin
           result_r_ns[630] = out_r[23:8];
           result_i_ns[630] = out_i[23:8];
        end
        10'd954 : begin
           result_r_ns[374] = out_r[23:8];
           result_i_ns[374] = out_i[23:8];
        end
        10'd955 : begin
           result_r_ns[886] = out_r[23:8];
           result_i_ns[886] = out_i[23:8];
        end
        10'd956 : begin
           result_r_ns[246] = out_r[23:8];
           result_i_ns[246] = out_i[23:8];
        end
        10'd957 : begin
           result_r_ns[758] = out_r[23:8];
           result_i_ns[758] = out_i[23:8];
        end
        10'd958 : begin
           result_r_ns[502] = out_r[23:8];
           result_i_ns[502] = out_i[23:8];
        end
        10'd959 : begin
           result_r_ns[1014] = out_r[23:8];
           result_i_ns[1014] = out_i[23:8];
        end
        10'd960 : begin
           result_r_ns[14] = out_r[23:8];
           result_i_ns[14] = out_i[23:8];
        end
        10'd961 : begin
           result_r_ns[526] = out_r[23:8];
           result_i_ns[526] = out_i[23:8];
        end
        10'd962 : begin
           result_r_ns[270] = out_r[23:8];
           result_i_ns[270] = out_i[23:8];
        end
        10'd963 : begin
           result_r_ns[782] = out_r[23:8];
           result_i_ns[782] = out_i[23:8];
        end
        10'd964 : begin
           result_r_ns[142] = out_r[23:8];
           result_i_ns[142] = out_i[23:8];
        end
        10'd965 : begin
           result_r_ns[654] = out_r[23:8];
           result_i_ns[654] = out_i[23:8];
        end
        10'd966 : begin
           result_r_ns[398] = out_r[23:8];
           result_i_ns[398] = out_i[23:8];
        end
        10'd967 : begin
           result_r_ns[910] = out_r[23:8];
           result_i_ns[910] = out_i[23:8];
        end
        10'd968 : begin
           result_r_ns[78] = out_r[23:8];
           result_i_ns[78] = out_i[23:8];
        end
        10'd969 : begin
           result_r_ns[590] = out_r[23:8];
           result_i_ns[590] = out_i[23:8];
        end
        10'd970 : begin
           result_r_ns[334] = out_r[23:8];
           result_i_ns[334] = out_i[23:8];
        end
        10'd971 : begin
           result_r_ns[846] = out_r[23:8];
           result_i_ns[846] = out_i[23:8];
        end
        10'd972 : begin
           result_r_ns[206] = out_r[23:8];
           result_i_ns[206] = out_i[23:8];
        end
        10'd973 : begin
           result_r_ns[718] = out_r[23:8];
           result_i_ns[718] = out_i[23:8];
        end
        10'd974 : begin
           result_r_ns[462] = out_r[23:8];
           result_i_ns[462] = out_i[23:8];
        end
        10'd975 : begin
           result_r_ns[974] = out_r[23:8];
           result_i_ns[974] = out_i[23:8];
        end
        10'd976 : begin
           result_r_ns[46] = out_r[23:8];
           result_i_ns[46] = out_i[23:8];
        end
        10'd977 : begin
           result_r_ns[558] = out_r[23:8];
           result_i_ns[558] = out_i[23:8];
        end
        10'd978 : begin
           result_r_ns[302] = out_r[23:8];
           result_i_ns[302] = out_i[23:8];
        end
        10'd979 : begin
           result_r_ns[814] = out_r[23:8];
           result_i_ns[814] = out_i[23:8];
        end
        10'd980 : begin
           result_r_ns[174] = out_r[23:8];
           result_i_ns[174] = out_i[23:8];
        end
        10'd981 : begin
           result_r_ns[686] = out_r[23:8];
           result_i_ns[686] = out_i[23:8];
        end
        10'd982 : begin
           result_r_ns[430] = out_r[23:8];
           result_i_ns[430] = out_i[23:8];
        end
        10'd983 : begin
           result_r_ns[942] = out_r[23:8];
           result_i_ns[942] = out_i[23:8];
        end
        10'd984 : begin
           result_r_ns[110] = out_r[23:8];
           result_i_ns[110] = out_i[23:8];
        end
        10'd985 : begin
           result_r_ns[622] = out_r[23:8];
           result_i_ns[622] = out_i[23:8];
        end
        10'd986 : begin
           result_r_ns[366] = out_r[23:8];
           result_i_ns[366] = out_i[23:8];
        end
        10'd987 : begin
           result_r_ns[878] = out_r[23:8];
           result_i_ns[878] = out_i[23:8];
        end
        10'd988 : begin
           result_r_ns[238] = out_r[23:8];
           result_i_ns[238] = out_i[23:8];
        end
        10'd989 : begin
           result_r_ns[750] = out_r[23:8];
           result_i_ns[750] = out_i[23:8];
        end
        10'd990 : begin
           result_r_ns[494] = out_r[23:8];
           result_i_ns[494] = out_i[23:8];
        end
        10'd991 : begin
           result_r_ns[1006] = out_r[23:8];
           result_i_ns[1006] = out_i[23:8];
        end
        10'd992 : begin
           result_r_ns[30] = out_r[23:8];
           result_i_ns[30] = out_i[23:8];
        end
        10'd993 : begin
           result_r_ns[542] = out_r[23:8];
           result_i_ns[542] = out_i[23:8];
        end
        10'd994 : begin
           result_r_ns[286] = out_r[23:8];
           result_i_ns[286] = out_i[23:8];
        end
        10'd995 : begin
           result_r_ns[798] = out_r[23:8];
           result_i_ns[798] = out_i[23:8];
        end
        10'd996 : begin
           result_r_ns[158] = out_r[23:8];
           result_i_ns[158] = out_i[23:8];
        end
        10'd997 : begin
           result_r_ns[670] = out_r[23:8];
           result_i_ns[670] = out_i[23:8];
        end
        10'd998 : begin
           result_r_ns[414] = out_r[23:8];
           result_i_ns[414] = out_i[23:8];
        end
        10'd999 : begin
           result_r_ns[926] = out_r[23:8];
           result_i_ns[926] = out_i[23:8];
        end
        10'd1000 : begin
           result_r_ns[94] = out_r[23:8];
           result_i_ns[94] = out_i[23:8];
        end
        10'd1001 : begin
           result_r_ns[606] = out_r[23:8];
           result_i_ns[606] = out_i[23:8];
        end
        10'd1002 : begin
           result_r_ns[350] = out_r[23:8];
           result_i_ns[350] = out_i[23:8];
        end
        10'd1003 : begin
           result_r_ns[862] = out_r[23:8];
           result_i_ns[862] = out_i[23:8];
        end
        10'd1004 : begin
           result_r_ns[222] = out_r[23:8];
           result_i_ns[222] = out_i[23:8];
        end
        10'd1005 : begin
           result_r_ns[734] = out_r[23:8];
           result_i_ns[734] = out_i[23:8];
        end
        10'd1006 : begin
           result_r_ns[478] = out_r[23:8];
           result_i_ns[478] = out_i[23:8];
        end
        10'd1007 : begin
           result_r_ns[990] = out_r[23:8];
           result_i_ns[990] = out_i[23:8];
        end
        10'd1008 : begin
           result_r_ns[62] = out_r[23:8];
           result_i_ns[62] = out_i[23:8];
        end
        10'd1009 : begin
           result_r_ns[574] = out_r[23:8];
           result_i_ns[574] = out_i[23:8];
        end
        10'd1010 : begin
           result_r_ns[318] = out_r[23:8];
           result_i_ns[318] = out_i[23:8];
        end
        10'd1011 : begin
           result_r_ns[830] = out_r[23:8];
           result_i_ns[830] = out_i[23:8];
        end
        10'd1012 : begin
           result_r_ns[190] = out_r[23:8];
           result_i_ns[190] = out_i[23:8];
        end
        10'd1013 : begin
           result_r_ns[702] = out_r[23:8];
           result_i_ns[702] = out_i[23:8];
        end
        10'd1014 : begin
           result_r_ns[446] = out_r[23:8];
           result_i_ns[446] = out_i[23:8];
        end
        10'd1015 : begin
           result_r_ns[958] = out_r[23:8];
           result_i_ns[958] = out_i[23:8];
        end
        10'd1016 : begin
           result_r_ns[126] = out_r[23:8];
           result_i_ns[126] = out_i[23:8];
        end
        10'd1017 : begin
           result_r_ns[638] = out_r[23:8];
           result_i_ns[638] = out_i[23:8];
        end
        10'd1018 : begin
           result_r_ns[382] = out_r[23:8];
           result_i_ns[382] = out_i[23:8];
        end
        10'd1019 : begin
           result_r_ns[894] = out_r[23:8];
           result_i_ns[894] = out_i[23:8];
        end
        10'd1020 : begin
           result_r_ns[254] = out_r[23:8];
           result_i_ns[254] = out_i[23:8];
        end
        10'd1021 : begin
           result_r_ns[766] = out_r[23:8];
           result_i_ns[766] = out_i[23:8];
        end
        10'd1022 : begin
           result_r_ns[510] = out_r[23:8];
           result_i_ns[510] = out_i[23:8];
        end
        10'd1023 : begin
           result_r_ns[1022] = out_r[23:8];
           result_i_ns[1022] = out_i[23:8];
           next_over = 1'b1; 
        end
        endcase
    end
end

endmodule
