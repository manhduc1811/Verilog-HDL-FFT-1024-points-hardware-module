module tb_FFT;

	parameter 					FFT_size		= 1024;
	parameter 					IN_width		= 12;
	parameter 					OUT_width		= 16;
	parameter 					latency_limit	= 2052;

	parameter 					cycle			= 10.0;
	
	integer 					j, latency;
    reg signed	[IN_width-1:0] int_r [0:FFT_size-1];
    reg signed	[IN_width-1:0] int_i [0:FFT_size-1];
	reg 						clk, rst_n, in_valid;
	wire 						out_valid;
	reg signed [IN_width-1:0] 	din_r, din_i;
	wire signed [OUT_width-1:0] dout_r, dout_i;

	always #(cycle/2.0) 
		clk = ~clk;

	FFT uut_FFT(
		.clk(clk),
		.rst_n(rst_n),
		.in_valid(in_valid),
		.din_r(din_r),
		.din_i(din_i),
		.out_valid(out_valid),
		.dout_r(dout_r),
		.dout_i(dout_i)
	);
	
	initial begin
		int_r[0] =  0;
		int_r[1] =  99;
		int_r[2] =  191;
		int_r[3] =  271;
		int_r[4] =  332;
		int_r[5] =  370;
		int_r[6] =  384;
		int_r[7] =  370;
		int_r[8] =  332;
		int_r[9] =  271;
		int_r[10] =  192;
		int_r[11] =  99;
		int_r[12] =  0;
		int_r[13] =  -100;
		int_r[14] =  -192;
		int_r[15] =  -272;
		int_r[16] =  -333;
		int_r[17] =  -371;
		int_r[18] =  -384;
		int_r[19] =  -371;
		int_r[20] =  -333;
		int_r[21] =  -272;
		int_r[22] =  -193;
		int_r[23] =  -100;
		int_r[24] =  -1;
		int_r[25] =  99;
		int_r[26] =  191;
		int_r[27] =  271;
		int_r[28] =  332;
		int_r[29] =  370;
		int_r[30] =  384;
		int_r[31] =  370;
		int_r[32] =  332;
		int_r[33] =  271;
		int_r[34] =  192;
		int_r[35] =  99;
		int_r[36] =  0;
		int_r[37] =  -100;
		int_r[38] =  -192;
		int_r[39] =  -272;
		int_r[40] =  -333;
		int_r[41] =  -371;
		int_r[42] =  -384;
		int_r[43] =  -371;
		int_r[44] =  -333;
		int_r[45] =  -272;
		int_r[46] =  -193;
		int_r[47] =  -100;
		int_r[48] =  -1;
		int_r[49] =  99;
		int_r[50] =  191;
		int_r[51] =  271;
		int_r[52] =  332;
		int_r[53] =  370;
		int_r[54] =  384;
		int_r[55] =  370;
		int_r[56] =  332;
		int_r[57] =  271;
		int_r[58] =  192;
		int_r[59] =  99;
		int_r[60] =  0;
		int_r[61] =  -100;
		int_r[62] =  -192;
		int_r[63] =  -272;
		int_r[64] =  -333;
		int_r[65] =  -371;
		int_r[66] =  -384;
		int_r[67] =  -371;
		int_r[68] =  -333;
		int_r[69] =  -272;
		int_r[70] =  -193;
		int_r[71] =  -100;
		int_r[72] =  -1;
		int_r[73] =  99;
		int_r[74] =  191;
		int_r[75] =  271;
		int_r[76] =  332;
		int_r[77] =  370;
		int_r[78] =  384;
		int_r[79] =  370;
		int_r[80] =  332;
		int_r[81] =  271;
		int_r[82] =  192;
		int_r[83] =  99;
		int_r[84] =  0;
		int_r[85] =  -100;
		int_r[86] =  -192;
		int_r[87] =  -272;
		int_r[88] =  -333;
		int_r[89] =  -371;
		int_r[90] =  -384;
		int_r[91] =  -371;
		int_r[92] =  -333;
		int_r[93] =  -272;
		int_r[94] =  -193;
		int_r[95] =  -100;
		int_r[96] =  -1;
		int_r[97] =  99;
		int_r[98] =  191;
		int_r[99] =  271;
		int_r[100] =  332;
		int_r[101] =  370;
		int_r[102] =  384;
		int_r[103] =  370;
		int_r[104] =  332;
		int_r[105] =  271;
		int_r[106] =  192;
		int_r[107] =  99;
		int_r[108] =  0;
		int_r[109] =  -100;
		int_r[110] =  -192;
		int_r[111] =  -272;
		int_r[112] =  -333;
		int_r[113] =  -371;
		int_r[114] =  -384;
		int_r[115] =  -371;
		int_r[116] =  -333;
		int_r[117] =  -272;
		int_r[118] =  -193;
		int_r[119] =  -100;
		int_r[120] =  -1;
		int_r[121] =  99;
		int_r[122] =  191;
		int_r[123] =  271;
		int_r[124] =  332;
		int_r[125] =  370;
		int_r[126] =  384;
		int_r[127] =  370;
		int_r[128] =  332;
		int_r[129] =  271;
		int_r[130] =  192;
		int_r[131] =  99;
		int_r[132] =  0;
		int_r[133] =  -100;
		int_r[134] =  -192;
		int_r[135] =  -272;
		int_r[136] =  -333;
		int_r[137] =  -371;
		int_r[138] =  -384;
		int_r[139] =  -371;
		int_r[140] =  -333;
		int_r[141] =  -272;
		int_r[142] =  -193;
		int_r[143] =  -100;
		int_r[144] =  -1;
		int_r[145] =  99;
		int_r[146] =  191;
		int_r[147] =  271;
		int_r[148] =  332;
		int_r[149] =  370;
		int_r[150] =  384;
		int_r[151] =  370;
		int_r[152] =  332;
		int_r[153] =  271;
		int_r[154] =  192;
		int_r[155] =  99;
		int_r[156] =  0;
		int_r[157] =  -100;
		int_r[158] =  -192;
		int_r[159] =  -272;
		int_r[160] =  -333;
		int_r[161] =  -371;
		int_r[162] =  -384;
		int_r[163] =  -371;
		int_r[164] =  -333;
		int_r[165] =  -272;
		int_r[166] =  -193;
		int_r[167] =  -100;
		int_r[168] =  -1;
		int_r[169] =  99;
		int_r[170] =  191;
		int_r[171] =  271;
		int_r[172] =  332;
		int_r[173] =  370;
		int_r[174] =  384;
		int_r[175] =  370;
		int_r[176] =  332;
		int_r[177] =  271;
		int_r[178] =  192;
		int_r[179] =  99;
		int_r[180] =  0;
		int_r[181] =  -100;
		int_r[182] =  -192;
		int_r[183] =  -272;
		int_r[184] =  -333;
		int_r[185] =  -371;
		int_r[186] =  -384;
		int_r[187] =  -371;
		int_r[188] =  -333;
		int_r[189] =  -272;
		int_r[190] =  -193;
		int_r[191] =  -100;
		int_r[192] =  -1;
		int_r[193] =  99;
		int_r[194] =  191;
		int_r[195] =  271;
		int_r[196] =  332;
		int_r[197] =  370;
		int_r[198] =  384;
		int_r[199] =  370;
		int_r[200] =  332;
		int_r[201] =  271;
		int_r[202] =  192;
		int_r[203] =  99;
		int_r[204] =  0;
		int_r[205] =  -100;
		int_r[206] =  -192;
		int_r[207] =  -272;
		int_r[208] =  -333;
		int_r[209] =  -371;
		int_r[210] =  -384;
		int_r[211] =  -371;
		int_r[212] =  -333;
		int_r[213] =  -272;
		int_r[214] =  -193;
		int_r[215] =  -100;
		int_r[216] =  -1;
		int_r[217] =  99;
		int_r[218] =  191;
		int_r[219] =  271;
		int_r[220] =  332;
		int_r[221] =  370;
		int_r[222] =  384;
		int_r[223] =  370;
		int_r[224] =  332;
		int_r[225] =  271;
		int_r[226] =  192;
		int_r[227] =  99;
		int_r[228] =  0;
		int_r[229] =  -100;
		int_r[230] =  -192;
		int_r[231] =  -272;
		int_r[232] =  -333;
		int_r[233] =  -371;
		int_r[234] =  -384;
		int_r[235] =  -371;
		int_r[236] =  -333;
		int_r[237] =  -272;
		int_r[238] =  -193;
		int_r[239] =  -100;
		int_r[240] =  -1;
		int_r[241] =  99;
		int_r[242] =  191;
		int_r[243] =  271;
		int_r[244] =  332;
		int_r[245] =  370;
		int_r[246] =  384;
		int_r[247] =  370;
		int_r[248] =  332;
		int_r[249] =  271;
		int_r[250] =  192;
		int_r[251] =  99;
		int_r[252] =  0;
		int_r[253] =  -100;
		int_r[254] =  -192;
		int_r[255] =  -272;
		int_r[256] =  -333;
		int_r[257] =  -371;
		int_r[258] =  -384;
		int_r[259] =  -371;
		int_r[260] =  -333;
		int_r[261] =  -272;
		int_r[262] =  -193;
		int_r[263] =  -100;
		int_r[264] =  -1;
		int_r[265] =  99;
		int_r[266] =  191;
		int_r[267] =  271;
		int_r[268] =  332;
		int_r[269] =  370;
		int_r[270] =  384;
		int_r[271] =  370;
		int_r[272] =  332;
		int_r[273] =  271;
		int_r[274] =  192;
		int_r[275] =  99;
		int_r[276] =  0;
		int_r[277] =  -100;
		int_r[278] =  -192;
		int_r[279] =  -272;
		int_r[280] =  -333;
		int_r[281] =  -371;
		int_r[282] =  -384;
		int_r[283] =  -371;
		int_r[284] =  -333;
		int_r[285] =  -272;
		int_r[286] =  -193;
		int_r[287] =  -100;
		int_r[288] =  -1;
		int_r[289] =  99;
		int_r[290] =  191;
		int_r[291] =  271;
		int_r[292] =  332;
		int_r[293] =  370;
		int_r[294] =  384;
		int_r[295] =  370;
		int_r[296] =  332;
		int_r[297] =  271;
		int_r[298] =  192;
		int_r[299] =  99;
		int_r[300] =  0;
		int_r[301] =  -100;
		int_r[302] =  -192;
		int_r[303] =  -272;
		int_r[304] =  -333;
		int_r[305] =  -371;
		int_r[306] =  -384;
		int_r[307] =  -371;
		int_r[308] =  -333;
		int_r[309] =  -272;
		int_r[310] =  -193;
		int_r[311] =  -100;
		int_r[312] =  -1;
		int_r[313] =  99;
		int_r[314] =  191;
		int_r[315] =  271;
		int_r[316] =  332;
		int_r[317] =  370;
		int_r[318] =  384;
		int_r[319] =  370;
		int_r[320] =  332;
		int_r[321] =  271;
		int_r[322] =  192;
		int_r[323] =  99;
		int_r[324] =  0;
		int_r[325] =  -100;
		int_r[326] =  -192;
		int_r[327] =  -272;
		int_r[328] =  -333;
		int_r[329] =  -371;
		int_r[330] =  -384;
		int_r[331] =  -371;
		int_r[332] =  -333;
		int_r[333] =  -272;
		int_r[334] =  -193;
		int_r[335] =  -100;
		int_r[336] =  -1;
		int_r[337] =  99;
		int_r[338] =  191;
		int_r[339] =  271;
		int_r[340] =  332;
		int_r[341] =  370;
		int_r[342] =  384;
		int_r[343] =  370;
		int_r[344] =  332;
		int_r[345] =  271;
		int_r[346] =  192;
		int_r[347] =  99;
		int_r[348] =  0;
		int_r[349] =  -100;
		int_r[350] =  -192;
		int_r[351] =  -272;
		int_r[352] =  -333;
		int_r[353] =  -371;
		int_r[354] =  -384;
		int_r[355] =  -371;
		int_r[356] =  -333;
		int_r[357] =  -272;
		int_r[358] =  -193;
		int_r[359] =  -100;
		int_r[360] =  -1;
		int_r[361] =  99;
		int_r[362] =  191;
		int_r[363] =  271;
		int_r[364] =  332;
		int_r[365] =  370;
		int_r[366] =  384;
		int_r[367] =  370;
		int_r[368] =  332;
		int_r[369] =  271;
		int_r[370] =  192;
		int_r[371] =  99;
		int_r[372] =  0;
		int_r[373] =  -100;
		int_r[374] =  -192;
		int_r[375] =  -272;
		int_r[376] =  -333;
		int_r[377] =  -371;
		int_r[378] =  -384;
		int_r[379] =  -371;
		int_r[380] =  -333;
		int_r[381] =  -272;
		int_r[382] =  -193;
		int_r[383] =  -100;
		int_r[384] =  -1;
		int_r[385] =  99;
		int_r[386] =  191;
		int_r[387] =  271;
		int_r[388] =  332;
		int_r[389] =  370;
		int_r[390] =  384;
		int_r[391] =  370;
		int_r[392] =  332;
		int_r[393] =  271;
		int_r[394] =  192;
		int_r[395] =  99;
		int_r[396] =  0;
		int_r[397] =  -100;
		int_r[398] =  -192;
		int_r[399] =  -272;
		int_r[400] =  -333;
		int_r[401] =  -371;
		int_r[402] =  -384;
		int_r[403] =  -371;
		int_r[404] =  -333;
		int_r[405] =  -272;
		int_r[406] =  -193;
		int_r[407] =  -100;
		int_r[408] =  -1;
		int_r[409] =  99;
		int_r[410] =  191;
		int_r[411] =  271;
		int_r[412] =  332;
		int_r[413] =  370;
		int_r[414] =  384;
		int_r[415] =  370;
		int_r[416] =  332;
		int_r[417] =  271;
		int_r[418] =  192;
		int_r[419] =  99;
		int_r[420] =  0;
		int_r[421] =  -100;
		int_r[422] =  -192;
		int_r[423] =  -272;
		int_r[424] =  -333;
		int_r[425] =  -371;
		int_r[426] =  -384;
		int_r[427] =  -371;
		int_r[428] =  -333;
		int_r[429] =  -272;
		int_r[430] =  -193;
		int_r[431] =  -100;
		int_r[432] =  -1;
		int_r[433] =  99;
		int_r[434] =  191;
		int_r[435] =  271;
		int_r[436] =  332;
		int_r[437] =  370;
		int_r[438] =  384;
		int_r[439] =  370;
		int_r[440] =  332;
		int_r[441] =  271;
		int_r[442] =  192;
		int_r[443] =  99;
		int_r[444] =  0;
		int_r[445] =  -100;
		int_r[446] =  -192;
		int_r[447] =  -272;
		int_r[448] =  -333;
		int_r[449] =  -371;
		int_r[450] =  -384;
		int_r[451] =  -371;
		int_r[452] =  -333;
		int_r[453] =  -272;
		int_r[454] =  -193;
		int_r[455] =  -100;
		int_r[456] =  -1;
		int_r[457] =  99;
		int_r[458] =  191;
		int_r[459] =  271;
		int_r[460] =  332;
		int_r[461] =  370;
		int_r[462] =  384;
		int_r[463] =  370;
		int_r[464] =  332;
		int_r[465] =  271;
		int_r[466] =  192;
		int_r[467] =  99;
		int_r[468] =  0;
		int_r[469] =  -100;
		int_r[470] =  -192;
		int_r[471] =  -272;
		int_r[472] =  -333;
		int_r[473] =  -371;
		int_r[474] =  -384;
		int_r[475] =  -371;
		int_r[476] =  -333;
		int_r[477] =  -272;
		int_r[478] =  -193;
		int_r[479] =  -100;
		int_r[480] =  -1;
		int_r[481] =  99;
		int_r[482] =  191;
		int_r[483] =  271;
		int_r[484] =  332;
		int_r[485] =  370;
		int_r[486] =  384;
		int_r[487] =  370;
		int_r[488] =  332;
		int_r[489] =  271;
		int_r[490] =  192;
		int_r[491] =  99;
		int_r[492] =  0;
		int_r[493] =  -100;
		int_r[494] =  -192;
		int_r[495] =  -272;
		int_r[496] =  -333;
		int_r[497] =  -371;
		int_r[498] =  -384;
		int_r[499] =  -371;
		int_r[500] =  -333;
		int_r[501] =  -272;
		int_r[502] =  -193;
		int_r[503] =  -100;
		int_r[504] =  -1;
		int_r[505] =  99;
		int_r[506] =  191;
		int_r[507] =  271;
		int_r[508] =  332;
		int_r[509] =  370;
		int_r[510] =  384;
		int_r[511] =  370;
		int_r[512] =  332;
		int_r[513] =  271;
		int_r[514] =  192;
		int_r[515] =  99;
		int_r[516] =  0;
		int_r[517] =  -100;
		int_r[518] =  -192;
		int_r[519] =  -272;
		int_r[520] =  -333;
		int_r[521] =  -371;
		int_r[522] =  -384;
		int_r[523] =  -371;
		int_r[524] =  -333;
		int_r[525] =  -272;
		int_r[526] =  -193;
		int_r[527] =  -100;
		int_r[528] =  -1;
		int_r[529] =  99;
		int_r[530] =  191;
		int_r[531] =  271;
		int_r[532] =  332;
		int_r[533] =  370;
		int_r[534] =  384;
		int_r[535] =  370;
		int_r[536] =  332;
		int_r[537] =  271;
		int_r[538] =  192;
		int_r[539] =  99;
		int_r[540] =  0;
		int_r[541] =  -100;
		int_r[542] =  -192;
		int_r[543] =  -272;
		int_r[544] =  -333;
		int_r[545] =  -371;
		int_r[546] =  -384;
		int_r[547] =  -371;
		int_r[548] =  -333;
		int_r[549] =  -272;
		int_r[550] =  -193;
		int_r[551] =  -100;
		int_r[552] =  -1;
		int_r[553] =  99;
		int_r[554] =  191;
		int_r[555] =  271;
		int_r[556] =  332;
		int_r[557] =  370;
		int_r[558] =  384;
		int_r[559] =  370;
		int_r[560] =  332;
		int_r[561] =  271;
		int_r[562] =  192;
		int_r[563] =  99;
		int_r[564] =  0;
		int_r[565] =  -100;
		int_r[566] =  -192;
		int_r[567] =  -272;
		int_r[568] =  -333;
		int_r[569] =  -371;
		int_r[570] =  -384;
		int_r[571] =  -371;
		int_r[572] =  -333;
		int_r[573] =  -272;
		int_r[574] =  -193;
		int_r[575] =  -100;
		int_r[576] =  -1;
		int_r[577] =  99;
		int_r[578] =  191;
		int_r[579] =  271;
		int_r[580] =  332;
		int_r[581] =  370;
		int_r[582] =  384;
		int_r[583] =  370;
		int_r[584] =  332;
		int_r[585] =  271;
		int_r[586] =  192;
		int_r[587] =  99;
		int_r[588] =  0;
		int_r[589] =  -100;
		int_r[590] =  -192;
		int_r[591] =  -272;
		int_r[592] =  -333;
		int_r[593] =  -371;
		int_r[594] =  -384;
		int_r[595] =  -371;
		int_r[596] =  -333;
		int_r[597] =  -272;
		int_r[598] =  -193;
		int_r[599] =  -100;
		int_r[600] =  -1;
		int_r[601] =  99;
		int_r[602] =  191;
		int_r[603] =  271;
		int_r[604] =  332;
		int_r[605] =  370;
		int_r[606] =  384;
		int_r[607] =  370;
		int_r[608] =  332;
		int_r[609] =  271;
		int_r[610] =  192;
		int_r[611] =  99;
		int_r[612] =  0;
		int_r[613] =  -100;
		int_r[614] =  -192;
		int_r[615] =  -272;
		int_r[616] =  -333;
		int_r[617] =  -371;
		int_r[618] =  -384;
		int_r[619] =  -371;
		int_r[620] =  -333;
		int_r[621] =  -272;
		int_r[622] =  -193;
		int_r[623] =  -100;
		int_r[624] =  -1;
		int_r[625] =  99;
		int_r[626] =  191;
		int_r[627] =  271;
		int_r[628] =  332;
		int_r[629] =  370;
		int_r[630] =  384;
		int_r[631] =  370;
		int_r[632] =  332;
		int_r[633] =  271;
		int_r[634] =  192;
		int_r[635] =  99;
		int_r[636] =  0;
		int_r[637] =  -100;
		int_r[638] =  -192;
		int_r[639] =  -272;
		int_r[640] =  -333;
		int_r[641] =  -371;
		int_r[642] =  -384;
		int_r[643] =  -371;
		int_r[644] =  -333;
		int_r[645] =  -272;
		int_r[646] =  -193;
		int_r[647] =  -100;
		int_r[648] =  -1;
		int_r[649] =  99;
		int_r[650] =  191;
		int_r[651] =  271;
		int_r[652] =  332;
		int_r[653] =  370;
		int_r[654] =  384;
		int_r[655] =  370;
		int_r[656] =  332;
		int_r[657] =  271;
		int_r[658] =  192;
		int_r[659] =  99;
		int_r[660] =  0;
		int_r[661] =  -100;
		int_r[662] =  -192;
		int_r[663] =  -272;
		int_r[664] =  -333;
		int_r[665] =  -371;
		int_r[666] =  -384;
		int_r[667] =  -371;
		int_r[668] =  -333;
		int_r[669] =  -272;
		int_r[670] =  -193;
		int_r[671] =  -100;
		int_r[672] =  -1;
		int_r[673] =  99;
		int_r[674] =  191;
		int_r[675] =  271;
		int_r[676] =  332;
		int_r[677] =  370;
		int_r[678] =  384;
		int_r[679] =  370;
		int_r[680] =  332;
		int_r[681] =  271;
		int_r[682] =  192;
		int_r[683] =  99;
		int_r[684] =  0;
		int_r[685] =  -100;
		int_r[686] =  -192;
		int_r[687] =  -272;
		int_r[688] =  -333;
		int_r[689] =  -371;
		int_r[690] =  -384;
		int_r[691] =  -371;
		int_r[692] =  -333;
		int_r[693] =  -272;
		int_r[694] =  -193;
		int_r[695] =  -100;
		int_r[696] =  -1;
		int_r[697] =  99;
		int_r[698] =  191;
		int_r[699] =  271;
		int_r[700] =  332;
		int_r[701] =  370;
		int_r[702] =  384;
		int_r[703] =  370;
		int_r[704] =  332;
		int_r[705] =  271;
		int_r[706] =  192;
		int_r[707] =  99;
		int_r[708] =  0;
		int_r[709] =  -100;
		int_r[710] =  -192;
		int_r[711] =  -272;
		int_r[712] =  -333;
		int_r[713] =  -371;
		int_r[714] =  -384;
		int_r[715] =  -371;
		int_r[716] =  -333;
		int_r[717] =  -272;
		int_r[718] =  -193;
		int_r[719] =  -100;
		int_r[720] =  -1;
		int_r[721] =  99;
		int_r[722] =  191;
		int_r[723] =  271;
		int_r[724] =  332;
		int_r[725] =  370;
		int_r[726] =  384;
		int_r[727] =  370;
		int_r[728] =  332;
		int_r[729] =  271;
		int_r[730] =  192;
		int_r[731] =  99;
		int_r[732] =  0;
		int_r[733] =  -100;
		int_r[734] =  -192;
		int_r[735] =  -272;
		int_r[736] =  -333;
		int_r[737] =  -371;
		int_r[738] =  -384;
		int_r[739] =  -371;
		int_r[740] =  -333;
		int_r[741] =  -272;
		int_r[742] =  -193;
		int_r[743] =  -100;
		int_r[744] =  -1;
		int_r[745] =  99;
		int_r[746] =  191;
		int_r[747] =  271;
		int_r[748] =  332;
		int_r[749] =  370;
		int_r[750] =  384;
		int_r[751] =  370;
		int_r[752] =  332;
		int_r[753] =  271;
		int_r[754] =  192;
		int_r[755] =  99;
		int_r[756] =  0;
		int_r[757] =  -100;
		int_r[758] =  -192;
		int_r[759] =  -272;
		int_r[760] =  -333;
		int_r[761] =  -371;
		int_r[762] =  -384;
		int_r[763] =  -371;
		int_r[764] =  -333;
		int_r[765] =  -272;
		int_r[766] =  -193;
		int_r[767] =  -100;
		int_r[768] =  -1;
		int_r[769] =  99;
		int_r[770] =  191;
		int_r[771] =  271;
		int_r[772] =  332;
		int_r[773] =  370;
		int_r[774] =  384;
		int_r[775] =  370;
		int_r[776] =  332;
		int_r[777] =  271;
		int_r[778] =  192;
		int_r[779] =  99;
		int_r[780] =  0;
		int_r[781] =  -100;
		int_r[782] =  -192;
		int_r[783] =  -272;
		int_r[784] =  -333;
		int_r[785] =  -371;
		int_r[786] =  -384;
		int_r[787] =  -371;
		int_r[788] =  -333;
		int_r[789] =  -272;
		int_r[790] =  -193;
		int_r[791] =  -100;
		int_r[792] =  -1;
		int_r[793] =  99;
		int_r[794] =  191;
		int_r[795] =  271;
		int_r[796] =  332;
		int_r[797] =  370;
		int_r[798] =  384;
		int_r[799] =  370;
		int_r[800] =  332;
		int_r[801] =  271;
		int_r[802] =  192;
		int_r[803] =  99;
		int_r[804] =  0;
		int_r[805] =  -100;
		int_r[806] =  -192;
		int_r[807] =  -272;
		int_r[808] =  -333;
		int_r[809] =  -371;
		int_r[810] =  -384;
		int_r[811] =  -371;
		int_r[812] =  -333;
		int_r[813] =  -272;
		int_r[814] =  -193;
		int_r[815] =  -100;
		int_r[816] =  -1;
		int_r[817] =  99;
		int_r[818] =  191;
		int_r[819] =  271;
		int_r[820] =  332;
		int_r[821] =  370;
		int_r[822] =  384;
		int_r[823] =  370;
		int_r[824] =  332;
		int_r[825] =  271;
		int_r[826] =  192;
		int_r[827] =  99;
		int_r[828] =  0;
		int_r[829] =  -100;
		int_r[830] =  -192;
		int_r[831] =  -272;
		int_r[832] =  -333;
		int_r[833] =  -371;
		int_r[834] =  -384;
		int_r[835] =  -371;
		int_r[836] =  -333;
		int_r[837] =  -272;
		int_r[838] =  -193;
		int_r[839] =  -100;
		int_r[840] =  -1;
		int_r[841] =  99;
		int_r[842] =  191;
		int_r[843] =  271;
		int_r[844] =  332;
		int_r[845] =  370;
		int_r[846] =  384;
		int_r[847] =  370;
		int_r[848] =  332;
		int_r[849] =  271;
		int_r[850] =  192;
		int_r[851] =  99;
		int_r[852] =  0;
		int_r[853] =  -100;
		int_r[854] =  -192;
		int_r[855] =  -272;
		int_r[856] =  -333;
		int_r[857] =  -371;
		int_r[858] =  -384;
		int_r[859] =  -371;
		int_r[860] =  -333;
		int_r[861] =  -272;
		int_r[862] =  -193;
		int_r[863] =  -100;
		int_r[864] =  -1;
		int_r[865] =  99;
		int_r[866] =  191;
		int_r[867] =  271;
		int_r[868] =  332;
		int_r[869] =  370;
		int_r[870] =  384;
		int_r[871] =  370;
		int_r[872] =  332;
		int_r[873] =  271;
		int_r[874] =  192;
		int_r[875] =  99;
		int_r[876] =  0;
		int_r[877] =  -100;
		int_r[878] =  -192;
		int_r[879] =  -272;
		int_r[880] =  -333;
		int_r[881] =  -371;
		int_r[882] =  -384;
		int_r[883] =  -371;
		int_r[884] =  -333;
		int_r[885] =  -272;
		int_r[886] =  -193;
		int_r[887] =  -100;
		int_r[888] =  -1;
		int_r[889] =  99;
		int_r[890] =  191;
		int_r[891] =  271;
		int_r[892] =  332;
		int_r[893] =  370;
		int_r[894] =  384;
		int_r[895] =  370;
		int_r[896] =  332;
		int_r[897] =  271;
		int_r[898] =  192;
		int_r[899] =  99;
		int_r[900] =  0;
		int_r[901] =  -100;
		int_r[902] =  -192;
		int_r[903] =  -272;
		int_r[904] =  -333;
		int_r[905] =  -371;
		int_r[906] =  -384;
		int_r[907] =  -371;
		int_r[908] =  -333;
		int_r[909] =  -272;
		int_r[910] =  -193;
		int_r[911] =  -100;
		int_r[912] =  -1;
		int_r[913] =  99;
		int_r[914] =  191;
		int_r[915] =  271;
		int_r[916] =  332;
		int_r[917] =  370;
		int_r[918] =  384;
		int_r[919] =  370;
		int_r[920] =  332;
		int_r[921] =  271;
		int_r[922] =  192;
		int_r[923] =  99;
		int_r[924] =  0;
		int_r[925] =  -100;
		int_r[926] =  -192;
		int_r[927] =  -272;
		int_r[928] =  -333;
		int_r[929] =  -371;
		int_r[930] =  -384;
		int_r[931] =  -371;
		int_r[932] =  -333;
		int_r[933] =  -272;
		int_r[934] =  -193;
		int_r[935] =  -100;
		int_r[936] =  -1;
		int_r[937] =  99;
		int_r[938] =  191;
		int_r[939] =  271;
		int_r[940] =  332;
		int_r[941] =  370;
		int_r[942] =  384;
		int_r[943] =  370;
		int_r[944] =  332;
		int_r[945] =  271;
		int_r[946] =  192;
		int_r[947] =  99;
		int_r[948] =  0;
		int_r[949] =  -100;
		int_r[950] =  -192;
		int_r[951] =  -272;
		int_r[952] =  -333;
		int_r[953] =  -371;
		int_r[954] =  -384;
		int_r[955] =  -371;
		int_r[956] =  -333;
		int_r[957] =  -272;
		int_r[958] =  -193;
		int_r[959] =  -100;
		int_r[960] =  -1;
		int_r[961] =  99;
		int_r[962] =  191;
		int_r[963] =  271;
		int_r[964] =  332;
		int_r[965] =  370;
		int_r[966] =  384;
		int_r[967] =  370;
		int_r[968] =  332;
		int_r[969] =  271;
		int_r[970] =  192;
		int_r[971] =  99;
		int_r[972] =  0;
		int_r[973] =  -100;
		int_r[974] =  -192;
		int_r[975] =  -272;
		int_r[976] =  -333;
		int_r[977] =  -371;
		int_r[978] =  -384;
		int_r[979] =  -371;
		int_r[980] =  -333;
		int_r[981] =  -272;
		int_r[982] =  -193;
		int_r[983] =  -100;
		int_r[984] =  -1;
		int_r[985] =  99;
		int_r[986] =  191;
		int_r[987] =  271;
		int_r[988] =  332;
		int_r[989] =  370;
		int_r[990] =  384;
		int_r[991] =  370;
		int_r[992] =  332;
		int_r[993] =  271;
		int_r[994] =  192;
		int_r[995] =  99;
		int_r[996] =  0;
		int_r[997] =  -100;
		int_r[998] =  -192;
		int_r[999] =  -272;
		int_r[1000] =  -333;
		int_r[1001] =  -371;
		int_r[1002] =  -384;
		int_r[1003] =  -371;
		int_r[1004] =  -333;
		int_r[1005] =  -272;
		int_r[1006] =  -193;
		int_r[1007] =  -100;
		int_r[1008] =  -1;
		int_r[1009] =  99;
		int_r[1010] =  191;
		int_r[1011] =  271;
		int_r[1012] =  332;
		int_r[1013] =  370;
		int_r[1014] =  384;
		int_r[1015] =  370;
		int_r[1016] =  332;
		int_r[1017] =  271;
		int_r[1018] =  192;
		int_r[1019] =  99;
		int_r[1020] =  0;
		int_r[1021] =  -100;
		int_r[1022] =  -192;
		int_r[1023] =  -272;
	end
	initial begin
		int_i[0] =    0;
		int_i[1] =    0;
		int_i[2] =    0;
		int_i[3] =    0;
		int_i[4] =    0;
		int_i[5] =    0;
		int_i[6] =    0;
		int_i[7] =    0;
		int_i[8] =    0;
		int_i[9] =    0;
		int_i[10] =    0;
		int_i[11] =    0;
		int_i[12] =    0;
		int_i[13] =    0;
		int_i[14] =    0;
		int_i[15] =    0;
		int_i[16] =    0;
		int_i[17] =    0;
		int_i[18] =    0;
		int_i[19] =    0;
		int_i[20] =    0;
		int_i[21] =    0;
		int_i[22] =    0;
		int_i[23] =    0;
		int_i[24] =    0;
		int_i[25] =    0;
		int_i[26] =    0;
		int_i[27] =    0;
		int_i[28] =    0;
		int_i[29] =    0;
		int_i[30] =    0;
		int_i[31] =    0;
		int_i[32] =    0;
		int_i[33] =    0;
		int_i[34] =    0;
		int_i[35] =    0;
		int_i[36] =    0;
		int_i[37] =    0;
		int_i[38] =    0;
		int_i[39] =    0;
		int_i[40] =    0;
		int_i[41] =    0;
		int_i[42] =    0;
		int_i[43] =    0;
		int_i[44] =    0;
		int_i[45] =    0;
		int_i[46] =    0;
		int_i[47] =    0;
		int_i[48] =    0;
		int_i[49] =    0;
		int_i[50] =    0;
		int_i[51] =    0;
		int_i[52] =    0;
		int_i[53] =    0;
		int_i[54] =    0;
		int_i[55] =    0;
		int_i[56] =    0;
		int_i[57] =    0;
		int_i[58] =    0;
		int_i[59] =    0;
		int_i[60] =    0;
		int_i[61] =    0;
		int_i[62] =    0;
		int_i[63] =    0;
		int_i[64] =    0;
		int_i[65] =    0;
		int_i[66] =    0;
		int_i[67] =    0;
		int_i[68] =    0;
		int_i[69] =    0;
		int_i[70] =    0;
		int_i[71] =    0;
		int_i[72] =    0;
		int_i[73] =    0;
		int_i[74] =    0;
		int_i[75] =    0;
		int_i[76] =    0;
		int_i[77] =    0;
		int_i[78] =    0;
		int_i[79] =    0;
		int_i[80] =    0;
		int_i[81] =    0;
		int_i[82] =    0;
		int_i[83] =    0;
		int_i[84] =    0;
		int_i[85] =    0;
		int_i[86] =    0;
		int_i[87] =    0;
		int_i[88] =    0;
		int_i[89] =    0;
		int_i[90] =    0;
		int_i[91] =    0;
		int_i[92] =    0;
		int_i[93] =    0;
		int_i[94] =    0;
		int_i[95] =    0;
		int_i[96] =    0;
		int_i[97] =    0;
		int_i[98] =    0;
		int_i[99] =    0;
		int_i[100] =    0;
		int_i[101] =    0;
		int_i[102] =    0;
		int_i[103] =    0;
		int_i[104] =    0;
		int_i[105] =    0;
		int_i[106] =    0;
		int_i[107] =    0;
		int_i[108] =    0;
		int_i[109] =    0;
		int_i[110] =    0;
		int_i[111] =    0;
		int_i[112] =    0;
		int_i[113] =    0;
		int_i[114] =    0;
		int_i[115] =    0;
		int_i[116] =    0;
		int_i[117] =    0;
		int_i[118] =    0;
		int_i[119] =    0;
		int_i[120] =    0;
		int_i[121] =    0;
		int_i[122] =    0;
		int_i[123] =    0;
		int_i[124] =    0;
		int_i[125] =    0;
		int_i[126] =    0;
		int_i[127] =    0;
		int_i[128] =    0;
		int_i[129] =    0;
		int_i[130] =    0;
		int_i[131] =    0;
		int_i[132] =    0;
		int_i[133] =    0;
		int_i[134] =    0;
		int_i[135] =    0;
		int_i[136] =    0;
		int_i[137] =    0;
		int_i[138] =    0;
		int_i[139] =    0;
		int_i[140] =    0;
		int_i[141] =    0;
		int_i[142] =    0;
		int_i[143] =    0;
		int_i[144] =    0;
		int_i[145] =    0;
		int_i[146] =    0;
		int_i[147] =    0;
		int_i[148] =    0;
		int_i[149] =    0;
		int_i[150] =    0;
		int_i[151] =    0;
		int_i[152] =    0;
		int_i[153] =    0;
		int_i[154] =    0;
		int_i[155] =    0;
		int_i[156] =    0;
		int_i[157] =    0;
		int_i[158] =    0;
		int_i[159] =    0;
		int_i[160] =    0;
		int_i[161] =    0;
		int_i[162] =    0;
		int_i[163] =    0;
		int_i[164] =    0;
		int_i[165] =    0;
		int_i[166] =    0;
		int_i[167] =    0;
		int_i[168] =    0;
		int_i[169] =    0;
		int_i[170] =    0;
		int_i[171] =    0;
		int_i[172] =    0;
		int_i[173] =    0;
		int_i[174] =    0;
		int_i[175] =    0;
		int_i[176] =    0;
		int_i[177] =    0;
		int_i[178] =    0;
		int_i[179] =    0;
		int_i[180] =    0;
		int_i[181] =    0;
		int_i[182] =    0;
		int_i[183] =    0;
		int_i[184] =    0;
		int_i[185] =    0;
		int_i[186] =    0;
		int_i[187] =    0;
		int_i[188] =    0;
		int_i[189] =    0;
		int_i[190] =    0;
		int_i[191] =    0;
		int_i[192] =    0;
		int_i[193] =    0;
		int_i[194] =    0;
		int_i[195] =    0;
		int_i[196] =    0;
		int_i[197] =    0;
		int_i[198] =    0;
		int_i[199] =    0;
		int_i[200] =    0;
		int_i[201] =    0;
		int_i[202] =    0;
		int_i[203] =    0;
		int_i[204] =    0;
		int_i[205] =    0;
		int_i[206] =    0;
		int_i[207] =    0;
		int_i[208] =    0;
		int_i[209] =    0;
		int_i[210] =    0;
		int_i[211] =    0;
		int_i[212] =    0;
		int_i[213] =    0;
		int_i[214] =    0;
		int_i[215] =    0;
		int_i[216] =    0;
		int_i[217] =    0;
		int_i[218] =    0;
		int_i[219] =    0;
		int_i[220] =    0;
		int_i[221] =    0;
		int_i[222] =    0;
		int_i[223] =    0;
		int_i[224] =    0;
		int_i[225] =    0;
		int_i[226] =    0;
		int_i[227] =    0;
		int_i[228] =    0;
		int_i[229] =    0;
		int_i[230] =    0;
		int_i[231] =    0;
		int_i[232] =    0;
		int_i[233] =    0;
		int_i[234] =    0;
		int_i[235] =    0;
		int_i[236] =    0;
		int_i[237] =    0;
		int_i[238] =    0;
		int_i[239] =    0;
		int_i[240] =    0;
		int_i[241] =    0;
		int_i[242] =    0;
		int_i[243] =    0;
		int_i[244] =    0;
		int_i[245] =    0;
		int_i[246] =    0;
		int_i[247] =    0;
		int_i[248] =    0;
		int_i[249] =    0;
		int_i[250] =    0;
		int_i[251] =    0;
		int_i[252] =    0;
		int_i[253] =    0;
		int_i[254] =    0;
		int_i[255] =    0;
		int_i[256] =    0;
		int_i[257] =    0;
		int_i[258] =    0;
		int_i[259] =    0;
		int_i[260] =    0;
		int_i[261] =    0;
		int_i[262] =    0;
		int_i[263] =    0;
		int_i[264] =    0;
		int_i[265] =    0;
		int_i[266] =    0;
		int_i[267] =    0;
		int_i[268] =    0;
		int_i[269] =    0;
		int_i[270] =    0;
		int_i[271] =    0;
		int_i[272] =    0;
		int_i[273] =    0;
		int_i[274] =    0;
		int_i[275] =    0;
		int_i[276] =    0;
		int_i[277] =    0;
		int_i[278] =    0;
		int_i[279] =    0;
		int_i[280] =    0;
		int_i[281] =    0;
		int_i[282] =    0;
		int_i[283] =    0;
		int_i[284] =    0;
		int_i[285] =    0;
		int_i[286] =    0;
		int_i[287] =    0;
		int_i[288] =    0;
		int_i[289] =    0;
		int_i[290] =    0;
		int_i[291] =    0;
		int_i[292] =    0;
		int_i[293] =    0;
		int_i[294] =    0;
		int_i[295] =    0;
		int_i[296] =    0;
		int_i[297] =    0;
		int_i[298] =    0;
		int_i[299] =    0;
		int_i[300] =    0;
		int_i[301] =    0;
		int_i[302] =    0;
		int_i[303] =    0;
		int_i[304] =    0;
		int_i[305] =    0;
		int_i[306] =    0;
		int_i[307] =    0;
		int_i[308] =    0;
		int_i[309] =    0;
		int_i[310] =    0;
		int_i[311] =    0;
		int_i[312] =    0;
		int_i[313] =    0;
		int_i[314] =    0;
		int_i[315] =    0;
		int_i[316] =    0;
		int_i[317] =    0;
		int_i[318] =    0;
		int_i[319] =    0;
		int_i[320] =    0;
		int_i[321] =    0;
		int_i[322] =    0;
		int_i[323] =    0;
		int_i[324] =    0;
		int_i[325] =    0;
		int_i[326] =    0;
		int_i[327] =    0;
		int_i[328] =    0;
		int_i[329] =    0;
		int_i[330] =    0;
		int_i[331] =    0;
		int_i[332] =    0;
		int_i[333] =    0;
		int_i[334] =    0;
		int_i[335] =    0;
		int_i[336] =    0;
		int_i[337] =    0;
		int_i[338] =    0;
		int_i[339] =    0;
		int_i[340] =    0;
		int_i[341] =    0;
		int_i[342] =    0;
		int_i[343] =    0;
		int_i[344] =    0;
		int_i[345] =    0;
		int_i[346] =    0;
		int_i[347] =    0;
		int_i[348] =    0;
		int_i[349] =    0;
		int_i[350] =    0;
		int_i[351] =    0;
		int_i[352] =    0;
		int_i[353] =    0;
		int_i[354] =    0;
		int_i[355] =    0;
		int_i[356] =    0;
		int_i[357] =    0;
		int_i[358] =    0;
		int_i[359] =    0;
		int_i[360] =    0;
		int_i[361] =    0;
		int_i[362] =    0;
		int_i[363] =    0;
		int_i[364] =    0;
		int_i[365] =    0;
		int_i[366] =    0;
		int_i[367] =    0;
		int_i[368] =    0;
		int_i[369] =    0;
		int_i[370] =    0;
		int_i[371] =    0;
		int_i[372] =    0;
		int_i[373] =    0;
		int_i[374] =    0;
		int_i[375] =    0;
		int_i[376] =    0;
		int_i[377] =    0;
		int_i[378] =    0;
		int_i[379] =    0;
		int_i[380] =    0;
		int_i[381] =    0;
		int_i[382] =    0;
		int_i[383] =    0;
		int_i[384] =    0;
		int_i[385] =    0;
		int_i[386] =    0;
		int_i[387] =    0;
		int_i[388] =    0;
		int_i[389] =    0;
		int_i[390] =    0;
		int_i[391] =    0;
		int_i[392] =    0;
		int_i[393] =    0;
		int_i[394] =    0;
		int_i[395] =    0;
		int_i[396] =    0;
		int_i[397] =    0;
		int_i[398] =    0;
		int_i[399] =    0;
		int_i[400] =    0;
		int_i[401] =    0;
		int_i[402] =    0;
		int_i[403] =    0;
		int_i[404] =    0;
		int_i[405] =    0;
		int_i[406] =    0;
		int_i[407] =    0;
		int_i[408] =    0;
		int_i[409] =    0;
		int_i[410] =    0;
		int_i[411] =    0;
		int_i[412] =    0;
		int_i[413] =    0;
		int_i[414] =    0;
		int_i[415] =    0;
		int_i[416] =    0;
		int_i[417] =    0;
		int_i[418] =    0;
		int_i[419] =    0;
		int_i[420] =    0;
		int_i[421] =    0;
		int_i[422] =    0;
		int_i[423] =    0;
		int_i[424] =    0;
		int_i[425] =    0;
		int_i[426] =    0;
		int_i[427] =    0;
		int_i[428] =    0;
		int_i[429] =    0;
		int_i[430] =    0;
		int_i[431] =    0;
		int_i[432] =    0;
		int_i[433] =    0;
		int_i[434] =    0;
		int_i[435] =    0;
		int_i[436] =    0;
		int_i[437] =    0;
		int_i[438] =    0;
		int_i[439] =    0;
		int_i[440] =    0;
		int_i[441] =    0;
		int_i[442] =    0;
		int_i[443] =    0;
		int_i[444] =    0;
		int_i[445] =    0;
		int_i[446] =    0;
		int_i[447] =    0;
		int_i[448] =    0;
		int_i[449] =    0;
		int_i[450] =    0;
		int_i[451] =    0;
		int_i[452] =    0;
		int_i[453] =    0;
		int_i[454] =    0;
		int_i[455] =    0;
		int_i[456] =    0;
		int_i[457] =    0;
		int_i[458] =    0;
		int_i[459] =    0;
		int_i[460] =    0;
		int_i[461] =    0;
		int_i[462] =    0;
		int_i[463] =    0;
		int_i[464] =    0;
		int_i[465] =    0;
		int_i[466] =    0;
		int_i[467] =    0;
		int_i[468] =    0;
		int_i[469] =    0;
		int_i[470] =    0;
		int_i[471] =    0;
		int_i[472] =    0;
		int_i[473] =    0;
		int_i[474] =    0;
		int_i[475] =    0;
		int_i[476] =    0;
		int_i[477] =    0;
		int_i[478] =    0;
		int_i[479] =    0;
		int_i[480] =    0;
		int_i[481] =    0;
		int_i[482] =    0;
		int_i[483] =    0;
		int_i[484] =    0;
		int_i[485] =    0;
		int_i[486] =    0;
		int_i[487] =    0;
		int_i[488] =    0;
		int_i[489] =    0;
		int_i[490] =    0;
		int_i[491] =    0;
		int_i[492] =    0;
		int_i[493] =    0;
		int_i[494] =    0;
		int_i[495] =    0;
		int_i[496] =    0;
		int_i[497] =    0;
		int_i[498] =    0;
		int_i[499] =    0;
		int_i[500] =    0;
		int_i[501] =    0;
		int_i[502] =    0;
		int_i[503] =    0;
		int_i[504] =    0;
		int_i[505] =    0;
		int_i[506] =    0;
		int_i[507] =    0;
		int_i[508] =    0;
		int_i[509] =    0;
		int_i[510] =    0;
		int_i[511] =    0;
		int_i[512] =    0;
		int_i[513] =    0;
		int_i[514] =    0;
		int_i[515] =    0;
		int_i[516] =    0;
		int_i[517] =    0;
		int_i[518] =    0;
		int_i[519] =    0;
		int_i[520] =    0;
		int_i[521] =    0;
		int_i[522] =    0;
		int_i[523] =    0;
		int_i[524] =    0;
		int_i[525] =    0;
		int_i[526] =    0;
		int_i[527] =    0;
		int_i[528] =    0;
		int_i[529] =    0;
		int_i[530] =    0;
		int_i[531] =    0;
		int_i[532] =    0;
		int_i[533] =    0;
		int_i[534] =    0;
		int_i[535] =    0;
		int_i[536] =    0;
		int_i[537] =    0;
		int_i[538] =    0;
		int_i[539] =    0;
		int_i[540] =    0;
		int_i[541] =    0;
		int_i[542] =    0;
		int_i[543] =    0;
		int_i[544] =    0;
		int_i[545] =    0;
		int_i[546] =    0;
		int_i[547] =    0;
		int_i[548] =    0;
		int_i[549] =    0;
		int_i[550] =    0;
		int_i[551] =    0;
		int_i[552] =    0;
		int_i[553] =    0;
		int_i[554] =    0;
		int_i[555] =    0;
		int_i[556] =    0;
		int_i[557] =    0;
		int_i[558] =    0;
		int_i[559] =    0;
		int_i[560] =    0;
		int_i[561] =    0;
		int_i[562] =    0;
		int_i[563] =    0;
		int_i[564] =    0;
		int_i[565] =    0;
		int_i[566] =    0;
		int_i[567] =    0;
		int_i[568] =    0;
		int_i[569] =    0;
		int_i[570] =    0;
		int_i[571] =    0;
		int_i[572] =    0;
		int_i[573] =    0;
		int_i[574] =    0;
		int_i[575] =    0;
		int_i[576] =    0;
		int_i[577] =    0;
		int_i[578] =    0;
		int_i[579] =    0;
		int_i[580] =    0;
		int_i[581] =    0;
		int_i[582] =    0;
		int_i[583] =    0;
		int_i[584] =    0;
		int_i[585] =    0;
		int_i[586] =    0;
		int_i[587] =    0;
		int_i[588] =    0;
		int_i[589] =    0;
		int_i[590] =    0;
		int_i[591] =    0;
		int_i[592] =    0;
		int_i[593] =    0;
		int_i[594] =    0;
		int_i[595] =    0;
		int_i[596] =    0;
		int_i[597] =    0;
		int_i[598] =    0;
		int_i[599] =    0;
		int_i[600] =    0;
		int_i[601] =    0;
		int_i[602] =    0;
		int_i[603] =    0;
		int_i[604] =    0;
		int_i[605] =    0;
		int_i[606] =    0;
		int_i[607] =    0;
		int_i[608] =    0;
		int_i[609] =    0;
		int_i[610] =    0;
		int_i[611] =    0;
		int_i[612] =    0;
		int_i[613] =    0;
		int_i[614] =    0;
		int_i[615] =    0;
		int_i[616] =    0;
		int_i[617] =    0;
		int_i[618] =    0;
		int_i[619] =    0;
		int_i[620] =    0;
		int_i[621] =    0;
		int_i[622] =    0;
		int_i[623] =    0;
		int_i[624] =    0;
		int_i[625] =    0;
		int_i[626] =    0;
		int_i[627] =    0;
		int_i[628] =    0;
		int_i[629] =    0;
		int_i[630] =    0;
		int_i[631] =    0;
		int_i[632] =    0;
		int_i[633] =    0;
		int_i[634] =    0;
		int_i[635] =    0;
		int_i[636] =    0;
		int_i[637] =    0;
		int_i[638] =    0;
		int_i[639] =    0;
		int_i[640] =    0;
		int_i[641] =    0;
		int_i[642] =    0;
		int_i[643] =    0;
		int_i[644] =    0;
		int_i[645] =    0;
		int_i[646] =    0;
		int_i[647] =    0;
		int_i[648] =    0;
		int_i[649] =    0;
		int_i[650] =    0;
		int_i[651] =    0;
		int_i[652] =    0;
		int_i[653] =    0;
		int_i[654] =    0;
		int_i[655] =    0;
		int_i[656] =    0;
		int_i[657] =    0;
		int_i[658] =    0;
		int_i[659] =    0;
		int_i[660] =    0;
		int_i[661] =    0;
		int_i[662] =    0;
		int_i[663] =    0;
		int_i[664] =    0;
		int_i[665] =    0;
		int_i[666] =    0;
		int_i[667] =    0;
		int_i[668] =    0;
		int_i[669] =    0;
		int_i[670] =    0;
		int_i[671] =    0;
		int_i[672] =    0;
		int_i[673] =    0;
		int_i[674] =    0;
		int_i[675] =    0;
		int_i[676] =    0;
		int_i[677] =    0;
		int_i[678] =    0;
		int_i[679] =    0;
		int_i[680] =    0;
		int_i[681] =    0;
		int_i[682] =    0;
		int_i[683] =    0;
		int_i[684] =    0;
		int_i[685] =    0;
		int_i[686] =    0;
		int_i[687] =    0;
		int_i[688] =    0;
		int_i[689] =    0;
		int_i[690] =    0;
		int_i[691] =    0;
		int_i[692] =    0;
		int_i[693] =    0;
		int_i[694] =    0;
		int_i[695] =    0;
		int_i[696] =    0;
		int_i[697] =    0;
		int_i[698] =    0;
		int_i[699] =    0;
		int_i[700] =    0;
		int_i[701] =    0;
		int_i[702] =    0;
		int_i[703] =    0;
		int_i[704] =    0;
		int_i[705] =    0;
		int_i[706] =    0;
		int_i[707] =    0;
		int_i[708] =    0;
		int_i[709] =    0;
		int_i[710] =    0;
		int_i[711] =    0;
		int_i[712] =    0;
		int_i[713] =    0;
		int_i[714] =    0;
		int_i[715] =    0;
		int_i[716] =    0;
		int_i[717] =    0;
		int_i[718] =    0;
		int_i[719] =    0;
		int_i[720] =    0;
		int_i[721] =    0;
		int_i[722] =    0;
		int_i[723] =    0;
		int_i[724] =    0;
		int_i[725] =    0;
		int_i[726] =    0;
		int_i[727] =    0;
		int_i[728] =    0;
		int_i[729] =    0;
		int_i[730] =    0;
		int_i[731] =    0;
		int_i[732] =    0;
		int_i[733] =    0;
		int_i[734] =    0;
		int_i[735] =    0;
		int_i[736] =    0;
		int_i[737] =    0;
		int_i[738] =    0;
		int_i[739] =    0;
		int_i[740] =    0;
		int_i[741] =    0;
		int_i[742] =    0;
		int_i[743] =    0;
		int_i[744] =    0;
		int_i[745] =    0;
		int_i[746] =    0;
		int_i[747] =    0;
		int_i[748] =    0;
		int_i[749] =    0;
		int_i[750] =    0;
		int_i[751] =    0;
		int_i[752] =    0;
		int_i[753] =    0;
		int_i[754] =    0;
		int_i[755] =    0;
		int_i[756] =    0;
		int_i[757] =    0;
		int_i[758] =    0;
		int_i[759] =    0;
		int_i[760] =    0;
		int_i[761] =    0;
		int_i[762] =    0;
		int_i[763] =    0;
		int_i[764] =    0;
		int_i[765] =    0;
		int_i[766] =    0;
		int_i[767] =    0;
		int_i[768] =    0;
		int_i[769] =    0;
		int_i[770] =    0;
		int_i[771] =    0;
		int_i[772] =    0;
		int_i[773] =    0;
		int_i[774] =    0;
		int_i[775] =    0;
		int_i[776] =    0;
		int_i[777] =    0;
		int_i[778] =    0;
		int_i[779] =    0;
		int_i[780] =    0;
		int_i[781] =    0;
		int_i[782] =    0;
		int_i[783] =    0;
		int_i[784] =    0;
		int_i[785] =    0;
		int_i[786] =    0;
		int_i[787] =    0;
		int_i[788] =    0;
		int_i[789] =    0;
		int_i[790] =    0;
		int_i[791] =    0;
		int_i[792] =    0;
		int_i[793] =    0;
		int_i[794] =    0;
		int_i[795] =    0;
		int_i[796] =    0;
		int_i[797] =    0;
		int_i[798] =    0;
		int_i[799] =    0;
		int_i[800] =    0;
		int_i[801] =    0;
		int_i[802] =    0;
		int_i[803] =    0;
		int_i[804] =    0;
		int_i[805] =    0;
		int_i[806] =    0;
		int_i[807] =    0;
		int_i[808] =    0;
		int_i[809] =    0;
		int_i[810] =    0;
		int_i[811] =    0;
		int_i[812] =    0;
		int_i[813] =    0;
		int_i[814] =    0;
		int_i[815] =    0;
		int_i[816] =    0;
		int_i[817] =    0;
		int_i[818] =    0;
		int_i[819] =    0;
		int_i[820] =    0;
		int_i[821] =    0;
		int_i[822] =    0;
		int_i[823] =    0;
		int_i[824] =    0;
		int_i[825] =    0;
		int_i[826] =    0;
		int_i[827] =    0;
		int_i[828] =    0;
		int_i[829] =    0;
		int_i[830] =    0;
		int_i[831] =    0;
		int_i[832] =    0;
		int_i[833] =    0;
		int_i[834] =    0;
		int_i[835] =    0;
		int_i[836] =    0;
		int_i[837] =    0;
		int_i[838] =    0;
		int_i[839] =    0;
		int_i[840] =    0;
		int_i[841] =    0;
		int_i[842] =    0;
		int_i[843] =    0;
		int_i[844] =    0;
		int_i[845] =    0;
		int_i[846] =    0;
		int_i[847] =    0;
		int_i[848] =    0;
		int_i[849] =    0;
		int_i[850] =    0;
		int_i[851] =    0;
		int_i[852] =    0;
		int_i[853] =    0;
		int_i[854] =    0;
		int_i[855] =    0;
		int_i[856] =    0;
		int_i[857] =    0;
		int_i[858] =    0;
		int_i[859] =    0;
		int_i[860] =    0;
		int_i[861] =    0;
		int_i[862] =    0;
		int_i[863] =    0;
		int_i[864] =    0;
		int_i[865] =    0;
		int_i[866] =    0;
		int_i[867] =    0;
		int_i[868] =    0;
		int_i[869] =    0;
		int_i[870] =    0;
		int_i[871] =    0;
		int_i[872] =    0;
		int_i[873] =    0;
		int_i[874] =    0;
		int_i[875] =    0;
		int_i[876] =    0;
		int_i[877] =    0;
		int_i[878] =    0;
		int_i[879] =    0;
		int_i[880] =    0;
		int_i[881] =    0;
		int_i[882] =    0;
		int_i[883] =    0;
		int_i[884] =    0;
		int_i[885] =    0;
		int_i[886] =    0;
		int_i[887] =    0;
		int_i[888] =    0;
		int_i[889] =    0;
		int_i[890] =    0;
		int_i[891] =    0;
		int_i[892] =    0;
		int_i[893] =    0;
		int_i[894] =    0;
		int_i[895] =    0;
		int_i[896] =    0;
		int_i[897] =    0;
		int_i[898] =    0;
		int_i[899] =    0;
		int_i[900] =    0;
		int_i[901] =    0;
		int_i[902] =    0;
		int_i[903] =    0;
		int_i[904] =    0;
		int_i[905] =    0;
		int_i[906] =    0;
		int_i[907] =    0;
		int_i[908] =    0;
		int_i[909] =    0;
		int_i[910] =    0;
		int_i[911] =    0;
		int_i[912] =    0;
		int_i[913] =    0;
		int_i[914] =    0;
		int_i[915] =    0;
		int_i[916] =    0;
		int_i[917] =    0;
		int_i[918] =    0;
		int_i[919] =    0;
		int_i[920] =    0;
		int_i[921] =    0;
		int_i[922] =    0;
		int_i[923] =    0;
		int_i[924] =    0;
		int_i[925] =    0;
		int_i[926] =    0;
		int_i[927] =    0;
		int_i[928] =    0;
		int_i[929] =    0;
		int_i[930] =    0;
		int_i[931] =    0;
		int_i[932] =    0;
		int_i[933] =    0;
		int_i[934] =    0;
		int_i[935] =    0;
		int_i[936] =    0;
		int_i[937] =    0;
		int_i[938] =    0;
		int_i[939] =    0;
		int_i[940] =    0;
		int_i[941] =    0;
		int_i[942] =    0;
		int_i[943] =    0;
		int_i[944] =    0;
		int_i[945] =    0;
		int_i[946] =    0;
		int_i[947] =    0;
		int_i[948] =    0;
		int_i[949] =    0;
		int_i[950] =    0;
		int_i[951] =    0;
		int_i[952] =    0;
		int_i[953] =    0;
		int_i[954] =    0;
		int_i[955] =    0;
		int_i[956] =    0;
		int_i[957] =    0;
		int_i[958] =    0;
		int_i[959] =    0;
		int_i[960] =    0;
		int_i[961] =    0;
		int_i[962] =    0;
		int_i[963] =    0;
		int_i[964] =    0;
		int_i[965] =    0;
		int_i[966] =    0;
		int_i[967] =    0;
		int_i[968] =    0;
		int_i[969] =    0;
		int_i[970] =    0;
		int_i[971] =    0;
		int_i[972] =    0;
		int_i[973] =    0;
		int_i[974] =    0;
		int_i[975] =    0;
		int_i[976] =    0;
		int_i[977] =    0;
		int_i[978] =    0;
		int_i[979] =    0;
		int_i[980] =    0;
		int_i[981] =    0;
		int_i[982] =    0;
		int_i[983] =    0;
		int_i[984] =    0;
		int_i[985] =    0;
		int_i[986] =    0;
		int_i[987] =    0;
		int_i[988] =    0;
		int_i[989] =    0;
		int_i[990] =    0;
		int_i[991] =    0;
		int_i[992] =    0;
		int_i[993] =    0;
		int_i[994] =    0;
		int_i[995] =    0;
		int_i[996] =    0;
		int_i[997] =    0;
		int_i[998] =    0;
		int_i[999] =    0;
		int_i[1000] =    0;
		int_i[1001] =    0;
		int_i[1002] =    0;
		int_i[1003] =    0;
		int_i[1004] =    0;
		int_i[1005] =    0;
		int_i[1006] =    0;
		int_i[1007] =    0;
		int_i[1008] =    0;
		int_i[1009] =    0;
		int_i[1010] =    0;
		int_i[1011] =    0;
		int_i[1012] =    0;
		int_i[1013] =    0;
		int_i[1014] =    0;
		int_i[1015] =    0;
		int_i[1016] =    0;
		int_i[1017] =    0;
		int_i[1018] =    0;
		int_i[1019] =    0;
		int_i[1020] =    0;
		int_i[1021] =    0;
		int_i[1022] =    0;
		int_i[1023] =    0;
	end
	
	initial begin
		clk = 0;
		rst_n = 1;
		in_valid = 0;

		@(negedge clk);
		@(negedge clk) 
			rst_n = 0;
		@(negedge clk) 
			rst_n = 1;
		@(negedge clk);

		for(j=0;j<FFT_size;j=j+1) 
		begin
			@(negedge clk);
			in_valid 	= 1;
			din_r 		= int_r[j];
			din_i 		= int_i[j];
		end
		@(negedge clk) 
			in_valid = 0;

		for(j=0;j<FFT_size;j=j+1) 
		begin
			while(!out_valid) 
			begin
				@(negedge clk) 
					latency = latency + 1;
				if(latency > latency_limit) 
				begin
					$display("Latency too long (> %0d cycles)", latency_limit);
					$stop;
				end
			end	
			@(negedge clk);
		end
		$stop;
	end
endmodule
	

