module FFT1024_tb;

	parameter 					FFT_size		= 1024;
	parameter 					IN_width		= 12;
	parameter 					OUT_width		= 16;
	parameter 					latency_limit	= 2052;

	parameter 					cycle			= 10.0;
	
	integer 					j;
    reg signed	[IN_width-1:0]  int_r           [0:FFT_size-1];
    reg signed	[IN_width-1:0]  int_i           [0:FFT_size-1];
	reg 						clk, rst_n, in_valid;
	wire 						out_valid;
	reg signed  [IN_width-1:0] 	din_r, din_i;
	wire signed [OUT_width-1:0] dout_r, dout_i;
////////////////////////////////////////////
	always #(cycle/2.0) 
		clk = ~clk;
////////////////////////////////////////////
	FFT1024 uut_FFT1024(
		.clk(clk),
		.rst_n(rst_n),
		.in_valid(in_valid),
		.din_r(din_r),
		.din_i(din_i),
		.out_valid(out_valid),
		.dout_r(dout_r),
		.dout_i(dout_i)
	);
////////////////////////////////////////////	
	initial begin
		int_r[0] =  0;
		int_r[1] =  331;
		int_r[2] =  229;
		int_r[3] =  -21;
		int_r[4] =  92;
		int_r[5] =  437;
		int_r[6] =  450;
		int_r[7] =  90;
		int_r[8] =  -93;
		int_r[9] =  119;
		int_r[10] =  256;
		int_r[11] =  -40;
		int_r[12] =  -394;
		int_r[13] =  -324;
		int_r[14] =  -37;
		int_r[15] =  -75;
		int_r[16] =  -394;
		int_r[17] =  -436;
		int_r[18] =  -72;
		int_r[19] =  173;
		int_r[20] =  0;
		int_r[21] =  -174;
		int_r[22] =  71;
		int_r[23] =  435;
		int_r[24] =  393;
		int_r[25] =  74;
		int_r[26] =  36;
		int_r[27] =  323;
		int_r[28] =  393;
		int_r[29] =  39;
		int_r[30] =  -256;
		int_r[31] =  -120;
		int_r[32] =  92;
		int_r[33] =  -91;
		int_r[34] =  -451;
		int_r[35] =  -438;
		int_r[36] =  -93;
		int_r[37] =  20;
		int_r[38] =  -230;
		int_r[39] =  -332;
		int_r[40] =  -1;
		int_r[41] =  331;
		int_r[42] =  229;
		int_r[43] =  -21;
		int_r[44] =  92;
		int_r[45] =  437;
		int_r[46] =  450;
		int_r[47] =  90;
		int_r[48] =  -93;
		int_r[49] =  119;
		int_r[50] =  256;
		int_r[51] =  -40;
		int_r[52] =  -394;
		int_r[53] =  -324;
		int_r[54] =  -37;
		int_r[55] =  -75;
		int_r[56] =  -394;
		int_r[57] =  -436;
		int_r[58] =  -72;
		int_r[59] =  173;
		int_r[60] =  0;
		int_r[61] =  -174;
		int_r[62] =  71;
		int_r[63] =  435;
		int_r[64] =  393;
		int_r[65] =  74;
		int_r[66] =  36;
		int_r[67] =  323;
		int_r[68] =  393;
		int_r[69] =  39;
		int_r[70] =  -256;
		int_r[71] =  -120;
		int_r[72] =  92;
		int_r[73] =  -91;
		int_r[74] =  -451;
		int_r[75] =  -438;
		int_r[76] =  -93;
		int_r[77] =  20;
		int_r[78] =  -230;
		int_r[79] =  -332;
		int_r[80] =  -1;
		int_r[81] =  331;
		int_r[82] =  229;
		int_r[83] =  -21;
		int_r[84] =  92;
		int_r[85] =  437;
		int_r[86] =  450;
		int_r[87] =  90;
		int_r[88] =  -93;
		int_r[89] =  119;
		int_r[90] =  256;
		int_r[91] =  -40;
		int_r[92] =  -394;
		int_r[93] =  -324;
		int_r[94] =  -37;
		int_r[95] =  -75;
		int_r[96] =  -394;
		int_r[97] =  -436;
		int_r[98] =  -72;
		int_r[99] =  173;
		int_r[100] =  0;
		int_r[101] =  -174;
		int_r[102] =  71;
		int_r[103] =  435;
		int_r[104] =  393;
		int_r[105] =  74;
		int_r[106] =  36;
		int_r[107] =  323;
		int_r[108] =  393;
		int_r[109] =  39;
		int_r[110] =  -256;
		int_r[111] =  -120;
		int_r[112] =  92;
		int_r[113] =  -91;
		int_r[114] =  -451;
		int_r[115] =  -438;
		int_r[116] =  -93;
		int_r[117] =  20;
		int_r[118] =  -230;
		int_r[119] =  -332;
		int_r[120] =  -1;
		int_r[121] =  331;
		int_r[122] =  229;
		int_r[123] =  -21;
		int_r[124] =  92;
		int_r[125] =  437;
		int_r[126] =  450;
		int_r[127] =  90;
		int_r[128] =  -93;
		int_r[129] =  119;
		int_r[130] =  255;
		int_r[131] =  -40;
		int_r[132] =  -394;
		int_r[133] =  -324;
		int_r[134] =  -37;
		int_r[135] =  -75;
		int_r[136] =  -394;
		int_r[137] =  -436;
		int_r[138] =  -72;
		int_r[139] =  173;
		int_r[140] =  -1;
		int_r[141] =  -174;
		int_r[142] =  71;
		int_r[143] =  435;
		int_r[144] =  393;
		int_r[145] =  74;
		int_r[146] =  36;
		int_r[147] =  323;
		int_r[148] =  393;
		int_r[149] =  39;
		int_r[150] =  -256;
		int_r[151] =  -120;
		int_r[152] =  92;
		int_r[153] =  -91;
		int_r[154] =  -451;
		int_r[155] =  -438;
		int_r[156] =  -93;
		int_r[157] =  20;
		int_r[158] =  -230;
		int_r[159] =  -332;
		int_r[160] =  -1;
		int_r[161] =  331;
		int_r[162] =  229;
		int_r[163] =  -21;
		int_r[164] =  92;
		int_r[165] =  437;
		int_r[166] =  450;
		int_r[167] =  90;
		int_r[168] =  -93;
		int_r[169] =  119;
		int_r[170] =  255;
		int_r[171] =  -40;
		int_r[172] =  -394;
		int_r[173] =  -324;
		int_r[174] =  -37;
		int_r[175] =  -75;
		int_r[176] =  -394;
		int_r[177] =  -436;
		int_r[178] =  -72;
		int_r[179] =  173;
		int_r[180] =  0;
		int_r[181] =  -174;
		int_r[182] =  71;
		int_r[183] =  435;
		int_r[184] =  393;
		int_r[185] =  74;
		int_r[186] =  36;
		int_r[187] =  323;
		int_r[188] =  393;
		int_r[189] =  39;
		int_r[190] =  -256;
		int_r[191] =  -120;
		int_r[192] =  92;
		int_r[193] =  -91;
		int_r[194] =  -451;
		int_r[195] =  -438;
		int_r[196] =  -93;
		int_r[197] =  20;
		int_r[198] =  -230;
		int_r[199] =  -332;
		int_r[200] =  -1;
		int_r[201] =  331;
		int_r[202] =  229;
		int_r[203] =  -21;
		int_r[204] =  92;
		int_r[205] =  437;
		int_r[206] =  450;
		int_r[207] =  90;
		int_r[208] =  -93;
		int_r[209] =  119;
		int_r[210] =  255;
		int_r[211] =  -40;
		int_r[212] =  -394;
		int_r[213] =  -324;
		int_r[214] =  -37;
		int_r[215] =  -75;
		int_r[216] =  -394;
		int_r[217] =  -436;
		int_r[218] =  -72;
		int_r[219] =  173;
		int_r[220] =  -1;
		int_r[221] =  -174;
		int_r[222] =  71;
		int_r[223] =  435;
		int_r[224] =  393;
		int_r[225] =  74;
		int_r[226] =  36;
		int_r[227] =  323;
		int_r[228] =  393;
		int_r[229] =  39;
		int_r[230] =  -256;
		int_r[231] =  -120;
		int_r[232] =  92;
		int_r[233] =  -91;
		int_r[234] =  -451;
		int_r[235] =  -438;
		int_r[236] =  -93;
		int_r[237] =  20;
		int_r[238] =  -230;
		int_r[239] =  -332;
		int_r[240] =  -1;
		int_r[241] =  331;
		int_r[242] =  229;
		int_r[243] =  -21;
		int_r[244] =  92;
		int_r[245] =  437;
		int_r[246] =  450;
		int_r[247] =  90;
		int_r[248] =  -93;
		int_r[249] =  119;
		int_r[250] =  255;
		int_r[251] =  -40;
		int_r[252] =  -394;
		int_r[253] =  -324;
		int_r[254] =  -37;
		int_r[255] =  -75;
		int_r[256] =  -394;
		int_r[257] =  -436;
		int_r[258] =  -72;
		int_r[259] =  173;
		int_r[260] =  0;
		int_r[261] =  -174;
		int_r[262] =  71;
		int_r[263] =  435;
		int_r[264] =  393;
		int_r[265] =  74;
		int_r[266] =  36;
		int_r[267] =  323;
		int_r[268] =  393;
		int_r[269] =  39;
		int_r[270] =  -256;
		int_r[271] =  -120;
		int_r[272] =  92;
		int_r[273] =  -91;
		int_r[274] =  -451;
		int_r[275] =  -438;
		int_r[276] =  -93;
		int_r[277] =  20;
		int_r[278] =  -230;
		int_r[279] =  -332;
		int_r[280] =  0;
		int_r[281] =  331;
		int_r[282] =  229;
		int_r[283] =  -21;
		int_r[284] =  92;
		int_r[285] =  437;
		int_r[286] =  450;
		int_r[287] =  90;
		int_r[288] =  -93;
		int_r[289] =  119;
		int_r[290] =  256;
		int_r[291] =  -40;
		int_r[292] =  -394;
		int_r[293] =  -324;
		int_r[294] =  -37;
		int_r[295] =  -75;
		int_r[296] =  -394;
		int_r[297] =  -436;
		int_r[298] =  -72;
		int_r[299] =  173;
		int_r[300] =  0;
		int_r[301] =  -174;
		int_r[302] =  71;
		int_r[303] =  435;
		int_r[304] =  393;
		int_r[305] =  74;
		int_r[306] =  36;
		int_r[307] =  323;
		int_r[308] =  393;
		int_r[309] =  39;
		int_r[310] =  -256;
		int_r[311] =  -120;
		int_r[312] =  92;
		int_r[313] =  -91;
		int_r[314] =  -451;
		int_r[315] =  -438;
		int_r[316] =  -93;
		int_r[317] =  20;
		int_r[318] =  -230;
		int_r[319] =  -332;
		int_r[320] =  -1;
		int_r[321] =  331;
		int_r[322] =  229;
		int_r[323] =  -21;
		int_r[324] =  92;
		int_r[325] =  437;
		int_r[326] =  450;
		int_r[327] =  90;
		int_r[328] =  -93;
		int_r[329] =  119;
		int_r[330] =  256;
		int_r[331] =  -40;
		int_r[332] =  -394;
		int_r[333] =  -324;
		int_r[334] =  -37;
		int_r[335] =  -75;
		int_r[336] =  -394;
		int_r[337] =  -436;
		int_r[338] =  -72;
		int_r[339] =  173;
		int_r[340] =  0;
		int_r[341] =  -174;
		int_r[342] =  71;
		int_r[343] =  435;
		int_r[344] =  393;
		int_r[345] =  74;
		int_r[346] =  36;
		int_r[347] =  323;
		int_r[348] =  393;
		int_r[349] =  39;
		int_r[350] =  -256;
		int_r[351] =  -120;
		int_r[352] =  92;
		int_r[353] =  -91;
		int_r[354] =  -451;
		int_r[355] =  -438;
		int_r[356] =  -93;
		int_r[357] =  20;
		int_r[358] =  -230;
		int_r[359] =  -332;
		int_r[360] =  -1;
		int_r[361] =  331;
		int_r[362] =  229;
		int_r[363] =  -21;
		int_r[364] =  92;
		int_r[365] =  437;
		int_r[366] =  450;
		int_r[367] =  90;
		int_r[368] =  -93;
		int_r[369] =  119;
		int_r[370] =  256;
		int_r[371] =  -40;
		int_r[372] =  -394;
		int_r[373] =  -324;
		int_r[374] =  -37;
		int_r[375] =  -75;
		int_r[376] =  -394;
		int_r[377] =  -436;
		int_r[378] =  -72;
		int_r[379] =  173;
		int_r[380] =  0;
		int_r[381] =  -174;
		int_r[382] =  71;
		int_r[383] =  435;
		int_r[384] =  393;
		int_r[385] =  74;
		int_r[386] =  36;
		int_r[387] =  323;
		int_r[388] =  393;
		int_r[389] =  39;
		int_r[390] =  -256;
		int_r[391] =  -120;
		int_r[392] =  92;
		int_r[393] =  -91;
		int_r[394] =  -451;
		int_r[395] =  -438;
		int_r[396] =  -93;
		int_r[397] =  20;
		int_r[398] =  -230;
		int_r[399] =  -332;
		int_r[400] =  -1;
		int_r[401] =  331;
		int_r[402] =  229;
		int_r[403] =  -21;
		int_r[404] =  92;
		int_r[405] =  437;
		int_r[406] =  450;
		int_r[407] =  90;
		int_r[408] =  -93;
		int_r[409] =  119;
		int_r[410] =  256;
		int_r[411] =  -40;
		int_r[412] =  -394;
		int_r[413] =  -324;
		int_r[414] =  -37;
		int_r[415] =  -75;
		int_r[416] =  -394;
		int_r[417] =  -436;
		int_r[418] =  -72;
		int_r[419] =  173;
		int_r[420] =  -1;
		int_r[421] =  -174;
		int_r[422] =  71;
		int_r[423] =  435;
		int_r[424] =  393;
		int_r[425] =  74;
		int_r[426] =  36;
		int_r[427] =  323;
		int_r[428] =  393;
		int_r[429] =  39;
		int_r[430] =  -256;
		int_r[431] =  -120;
		int_r[432] =  92;
		int_r[433] =  -91;
		int_r[434] =  -451;
		int_r[435] =  -438;
		int_r[436] =  -93;
		int_r[437] =  20;
		int_r[438] =  -230;
		int_r[439] =  -332;
		int_r[440] =  0;
		int_r[441] =  331;
		int_r[442] =  229;
		int_r[443] =  -21;
		int_r[444] =  92;
		int_r[445] =  437;
		int_r[446] =  450;
		int_r[447] =  90;
		int_r[448] =  -93;
		int_r[449] =  119;
		int_r[450] =  256;
		int_r[451] =  -40;
		int_r[452] =  -394;
		int_r[453] =  -324;
		int_r[454] =  -37;
		int_r[455] =  -75;
		int_r[456] =  -394;
		int_r[457] =  -436;
		int_r[458] =  -72;
		int_r[459] =  173;
		int_r[460] =  0;
		int_r[461] =  -174;
		int_r[462] =  71;
		int_r[463] =  435;
		int_r[464] =  393;
		int_r[465] =  74;
		int_r[466] =  36;
		int_r[467] =  323;
		int_r[468] =  393;
		int_r[469] =  39;
		int_r[470] =  -257;
		int_r[471] =  -120;
		int_r[472] =  92;
		int_r[473] =  -91;
		int_r[474] =  -451;
		int_r[475] =  -438;
		int_r[476] =  -93;
		int_r[477] =  20;
		int_r[478] =  -230;
		int_r[479] =  -332;
		int_r[480] =  -1;
		int_r[481] =  331;
		int_r[482] =  229;
		int_r[483] =  -21;
		int_r[484] =  92;
		int_r[485] =  437;
		int_r[486] =  450;
		int_r[487] =  90;
		int_r[488] =  -93;
		int_r[489] =  119;
		int_r[490] =  256;
		int_r[491] =  -40;
		int_r[492] =  -394;
		int_r[493] =  -324;
		int_r[494] =  -37;
		int_r[495] =  -75;
		int_r[496] =  -394;
		int_r[497] =  -436;
		int_r[498] =  -72;
		int_r[499] =  173;
		int_r[500] =  0;
		int_r[501] =  -174;
		int_r[502] =  71;
		int_r[503] =  435;
		int_r[504] =  393;
		int_r[505] =  74;
		int_r[506] =  36;
		int_r[507] =  323;
		int_r[508] =  393;
		int_r[509] =  39;
		int_r[510] =  -256;
		int_r[511] =  -120;
		int_r[512] =  92;
		int_r[513] =  -91;
		int_r[514] =  -451;
		int_r[515] =  -438;
		int_r[516] =  -93;
		int_r[517] =  20;
		int_r[518] =  -230;
		int_r[519] =  -332;
		int_r[520] =  -1;
		int_r[521] =  331;
		int_r[522] =  229;
		int_r[523] =  -21;
		int_r[524] =  92;
		int_r[525] =  437;
		int_r[526] =  450;
		int_r[527] =  90;
		int_r[528] =  -93;
		int_r[529] =  119;
		int_r[530] =  256;
		int_r[531] =  -40;
		int_r[532] =  -394;
		int_r[533] =  -324;
		int_r[534] =  -37;
		int_r[535] =  -75;
		int_r[536] =  -394;
		int_r[537] =  -436;
		int_r[538] =  -72;
		int_r[539] =  173;
		int_r[540] =  -1;
		int_r[541] =  -174;
		int_r[542] =  71;
		int_r[543] =  435;
		int_r[544] =  393;
		int_r[545] =  74;
		int_r[546] =  36;
		int_r[547] =  323;
		int_r[548] =  393;
		int_r[549] =  39;
		int_r[550] =  -257;
		int_r[551] =  -120;
		int_r[552] =  92;
		int_r[553] =  -91;
		int_r[554] =  -451;
		int_r[555] =  -438;
		int_r[556] =  -93;
		int_r[557] =  20;
		int_r[558] =  -230;
		int_r[559] =  -332;
		int_r[560] =  0;
		int_r[561] =  331;
		int_r[562] =  229;
		int_r[563] =  -21;
		int_r[564] =  92;
		int_r[565] =  437;
		int_r[566] =  450;
		int_r[567] =  90;
		int_r[568] =  -93;
		int_r[569] =  119;
		int_r[570] =  256;
		int_r[571] =  -40;
		int_r[572] =  -394;
		int_r[573] =  -324;
		int_r[574] =  -37;
		int_r[575] =  -75;
		int_r[576] =  -394;
		int_r[577] =  -436;
		int_r[578] =  -72;
		int_r[579] =  173;
		int_r[580] =  0;
		int_r[581] =  -174;
		int_r[582] =  71;
		int_r[583] =  435;
		int_r[584] =  393;
		int_r[585] =  74;
		int_r[586] =  36;
		int_r[587] =  323;
		int_r[588] =  393;
		int_r[589] =  39;
		int_r[590] =  -256;
		int_r[591] =  -120;
		int_r[592] =  92;
		int_r[593] =  -91;
		int_r[594] =  -451;
		int_r[595] =  -438;
		int_r[596] =  -93;
		int_r[597] =  20;
		int_r[598] =  -230;
		int_r[599] =  -332;
		int_r[600] =  -1;
		int_r[601] =  331;
		int_r[602] =  229;
		int_r[603] =  -21;
		int_r[604] =  92;
		int_r[605] =  437;
		int_r[606] =  450;
		int_r[607] =  90;
		int_r[608] =  -93;
		int_r[609] =  119;
		int_r[610] =  256;
		int_r[611] =  -40;
		int_r[612] =  -394;
		int_r[613] =  -324;
		int_r[614] =  -37;
		int_r[615] =  -75;
		int_r[616] =  -394;
		int_r[617] =  -436;
		int_r[618] =  -72;
		int_r[619] =  173;
		int_r[620] =  0;
		int_r[621] =  -174;
		int_r[622] =  71;
		int_r[623] =  435;
		int_r[624] =  393;
		int_r[625] =  74;
		int_r[626] =  36;
		int_r[627] =  323;
		int_r[628] =  393;
		int_r[629] =  39;
		int_r[630] =  -257;
		int_r[631] =  -120;
		int_r[632] =  92;
		int_r[633] =  -91;
		int_r[634] =  -451;
		int_r[635] =  -438;
		int_r[636] =  -93;
		int_r[637] =  20;
		int_r[638] =  -230;
		int_r[639] =  -332;
		int_r[640] =  -1;
		int_r[641] =  331;
		int_r[642] =  229;
		int_r[643] =  -21;
		int_r[644] =  92;
		int_r[645] =  437;
		int_r[646] =  450;
		int_r[647] =  90;
		int_r[648] =  -93;
		int_r[649] =  119;
		int_r[650] =  256;
		int_r[651] =  -40;
		int_r[652] =  -394;
		int_r[653] =  -324;
		int_r[654] =  -37;
		int_r[655] =  -75;
		int_r[656] =  -394;
		int_r[657] =  -436;
		int_r[658] =  -72;
		int_r[659] =  173;
		int_r[660] =  0;
		int_r[661] =  -174;
		int_r[662] =  71;
		int_r[663] =  435;
		int_r[664] =  393;
		int_r[665] =  74;
		int_r[666] =  36;
		int_r[667] =  323;
		int_r[668] =  393;
		int_r[669] =  39;
		int_r[670] =  -256;
		int_r[671] =  -120;
		int_r[672] =  92;
		int_r[673] =  -91;
		int_r[674] =  -451;
		int_r[675] =  -438;
		int_r[676] =  -93;
		int_r[677] =  20;
		int_r[678] =  -230;
		int_r[679] =  -332;
		int_r[680] =  0;
		int_r[681] =  331;
		int_r[682] =  229;
		int_r[683] =  -21;
		int_r[684] =  92;
		int_r[685] =  437;
		int_r[686] =  450;
		int_r[687] =  90;
		int_r[688] =  -93;
		int_r[689] =  119;
		int_r[690] =  256;
		int_r[691] =  -40;
		int_r[692] =  -394;
		int_r[693] =  -324;
		int_r[694] =  -37;
		int_r[695] =  -75;
		int_r[696] =  -394;
		int_r[697] =  -436;
		int_r[698] =  -72;
		int_r[699] =  173;
		int_r[700] =  -1;
		int_r[701] =  -174;
		int_r[702] =  71;
		int_r[703] =  435;
		int_r[704] =  393;
		int_r[705] =  74;
		int_r[706] =  36;
		int_r[707] =  323;
		int_r[708] =  393;
		int_r[709] =  39;
		int_r[710] =  -257;
		int_r[711] =  -120;
		int_r[712] =  92;
		int_r[713] =  -91;
		int_r[714] =  -451;
		int_r[715] =  -438;
		int_r[716] =  -93;
		int_r[717] =  20;
		int_r[718] =  -230;
		int_r[719] =  -332;
		int_r[720] =  -1;
		int_r[721] =  331;
		int_r[722] =  229;
		int_r[723] =  -21;
		int_r[724] =  92;
		int_r[725] =  437;
		int_r[726] =  450;
		int_r[727] =  90;
		int_r[728] =  -93;
		int_r[729] =  119;
		int_r[730] =  256;
		int_r[731] =  -40;
		int_r[732] =  -394;
		int_r[733] =  -324;
		int_r[734] =  -37;
		int_r[735] =  -75;
		int_r[736] =  -394;
		int_r[737] =  -436;
		int_r[738] =  -72;
		int_r[739] =  173;
		int_r[740] =  0;
		int_r[741] =  -174;
		int_r[742] =  71;
		int_r[743] =  435;
		int_r[744] =  393;
		int_r[745] =  74;
		int_r[746] =  36;
		int_r[747] =  323;
		int_r[748] =  393;
		int_r[749] =  39;
		int_r[750] =  -256;
		int_r[751] =  -120;
		int_r[752] =  92;
		int_r[753] =  -91;
		int_r[754] =  -451;
		int_r[755] =  -438;
		int_r[756] =  -93;
		int_r[757] =  20;
		int_r[758] =  -230;
		int_r[759] =  -332;
		int_r[760] =  -1;
		int_r[761] =  331;
		int_r[762] =  229;
		int_r[763] =  -21;
		int_r[764] =  92;
		int_r[765] =  437;
		int_r[766] =  450;
		int_r[767] =  90;
		int_r[768] =  -93;
		int_r[769] =  119;
		int_r[770] =  256;
		int_r[771] =  -40;
		int_r[772] =  -394;
		int_r[773] =  -324;
		int_r[774] =  -37;
		int_r[775] =  -75;
		int_r[776] =  -394;
		int_r[777] =  -436;
		int_r[778] =  -72;
		int_r[779] =  173;
		int_r[780] =  0;
		int_r[781] =  -174;
		int_r[782] =  71;
		int_r[783] =  435;
		int_r[784] =  393;
		int_r[785] =  74;
		int_r[786] =  36;
		int_r[787] =  323;
		int_r[788] =  393;
		int_r[789] =  39;
		int_r[790] =  -257;
		int_r[791] =  -120;
		int_r[792] =  92;
		int_r[793] =  -91;
		int_r[794] =  -451;
		int_r[795] =  -438;
		int_r[796] =  -93;
		int_r[797] =  20;
		int_r[798] =  -230;
		int_r[799] =  -332;
		int_r[800] =  -1;
		int_r[801] =  331;
		int_r[802] =  229;
		int_r[803] =  -21;
		int_r[804] =  92;
		int_r[805] =  437;
		int_r[806] =  450;
		int_r[807] =  90;
		int_r[808] =  -93;
		int_r[809] =  119;
		int_r[810] =  256;
		int_r[811] =  -40;
		int_r[812] =  -394;
		int_r[813] =  -324;
		int_r[814] =  -37;
		int_r[815] =  -75;
		int_r[816] =  -394;
		int_r[817] =  -436;
		int_r[818] =  -72;
		int_r[819] =  173;
		int_r[820] =  -1;
		int_r[821] =  -174;
		int_r[822] =  71;
		int_r[823] =  435;
		int_r[824] =  393;
		int_r[825] =  74;
		int_r[826] =  36;
		int_r[827] =  323;
		int_r[828] =  393;
		int_r[829] =  39;
		int_r[830] =  -257;
		int_r[831] =  -120;
		int_r[832] =  92;
		int_r[833] =  -91;
		int_r[834] =  -451;
		int_r[835] =  -438;
		int_r[836] =  -93;
		int_r[837] =  20;
		int_r[838] =  -230;
		int_r[839] =  -332;
		int_r[840] =  0;
		int_r[841] =  331;
		int_r[842] =  229;
		int_r[843] =  -21;
		int_r[844] =  92;
		int_r[845] =  437;
		int_r[846] =  450;
		int_r[847] =  90;
		int_r[848] =  -93;
		int_r[849] =  119;
		int_r[850] =  256;
		int_r[851] =  -40;
		int_r[852] =  -394;
		int_r[853] =  -324;
		int_r[854] =  -37;
		int_r[855] =  -75;
		int_r[856] =  -394;
		int_r[857] =  -436;
		int_r[858] =  -72;
		int_r[859] =  173;
		int_r[860] =  -1;
		int_r[861] =  -174;
		int_r[862] =  71;
		int_r[863] =  435;
		int_r[864] =  393;
		int_r[865] =  74;
		int_r[866] =  36;
		int_r[867] =  323;
		int_r[868] =  393;
		int_r[869] =  39;
		int_r[870] =  -256;
		int_r[871] =  -120;
		int_r[872] =  92;
		int_r[873] =  -91;
		int_r[874] =  -451;
		int_r[875] =  -438;
		int_r[876] =  -93;
		int_r[877] =  20;
		int_r[878] =  -230;
		int_r[879] =  -332;
		int_r[880] =  0;
		int_r[881] =  331;
		int_r[882] =  229;
		int_r[883] =  -21;
		int_r[884] =  92;
		int_r[885] =  437;
		int_r[886] =  450;
		int_r[887] =  90;
		int_r[888] =  -93;
		int_r[889] =  119;
		int_r[890] =  255;
		int_r[891] =  -40;
		int_r[892] =  -394;
		int_r[893] =  -324;
		int_r[894] =  -37;
		int_r[895] =  -75;
		int_r[896] =  -394;
		int_r[897] =  -436;
		int_r[898] =  -72;
		int_r[899] =  173;
		int_r[900] =  0;
		int_r[901] =  -174;
		int_r[902] =  71;
		int_r[903] =  435;
		int_r[904] =  393;
		int_r[905] =  74;
		int_r[906] =  36;
		int_r[907] =  323;
		int_r[908] =  393;
		int_r[909] =  39;
		int_r[910] =  -256;
		int_r[911] =  -120;
		int_r[912] =  92;
		int_r[913] =  -91;
		int_r[914] =  -451;
		int_r[915] =  -438;
		int_r[916] =  -93;
		int_r[917] =  20;
		int_r[918] =  -230;
		int_r[919] =  -332;
		int_r[920] =  -1;
		int_r[921] =  331;
		int_r[922] =  229;
		int_r[923] =  -21;
		int_r[924] =  92;
		int_r[925] =  437;
		int_r[926] =  450;
		int_r[927] =  90;
		int_r[928] =  -93;
		int_r[929] =  119;
		int_r[930] =  256;
		int_r[931] =  -40;
		int_r[932] =  -394;
		int_r[933] =  -324;
		int_r[934] =  -37;
		int_r[935] =  -75;
		int_r[936] =  -394;
		int_r[937] =  -436;
		int_r[938] =  -72;
		int_r[939] =  173;
		int_r[940] =  0;
		int_r[941] =  -174;
		int_r[942] =  71;
		int_r[943] =  435;
		int_r[944] =  393;
		int_r[945] =  74;
		int_r[946] =  36;
		int_r[947] =  323;
		int_r[948] =  393;
		int_r[949] =  39;
		int_r[950] =  -256;
		int_r[951] =  -120;
		int_r[952] =  92;
		int_r[953] =  -91;
		int_r[954] =  -451;
		int_r[955] =  -438;
		int_r[956] =  -93;
		int_r[957] =  20;
		int_r[958] =  -230;
		int_r[959] =  -332;
		int_r[960] =  -1;
		int_r[961] =  331;
		int_r[962] =  229;
		int_r[963] =  -21;
		int_r[964] =  92;
		int_r[965] =  437;
		int_r[966] =  450;
		int_r[967] =  90;
		int_r[968] =  -93;
		int_r[969] =  119;
		int_r[970] =  256;
		int_r[971] =  -40;
		int_r[972] =  -394;
		int_r[973] =  -324;
		int_r[974] =  -37;
		int_r[975] =  -75;
		int_r[976] =  -394;
		int_r[977] =  -436;
		int_r[978] =  -72;
		int_r[979] =  173;
		int_r[980] =  0;
		int_r[981] =  -174;
		int_r[982] =  71;
		int_r[983] =  435;
		int_r[984] =  393;
		int_r[985] =  74;
		int_r[986] =  36;
		int_r[987] =  323;
		int_r[988] =  393;
		int_r[989] =  39;
		int_r[990] =  -257;
		int_r[991] =  -120;
		int_r[992] =  92;
		int_r[993] =  -91;
		int_r[994] =  -451;
		int_r[995] =  -438;
		int_r[996] =  -93;
		int_r[997] =  20;
		int_r[998] =  -230;
		int_r[999] =  -332;
		int_r[1000] =  -1;
		int_r[1001] =  331;
		int_r[1002] =  229;
		int_r[1003] =  -21;
		int_r[1004] =  92;
		int_r[1005] =  437;
		int_r[1006] =  450;
		int_r[1007] =  90;
		int_r[1008] =  -93;
		int_r[1009] =  119;
		int_r[1010] =  256;
		int_r[1011] =  -40;
		int_r[1012] =  -394;
		int_r[1013] =  -324;
		int_r[1014] =  -37;
		int_r[1015] =  -75;
		int_r[1016] =  -394;
		int_r[1017] =  -436;
		int_r[1018] =  -72;
		int_r[1019] =  173;
		int_r[1020] =  0;
		int_r[1021] =  -174;
		int_r[1022] =  71;
		int_r[1023] =  435;
	end
	initial begin
		int_i[0] =  0;
		int_i[1] =  0;
		int_i[2] =  0;
		int_i[3] =  0;
		int_i[4] =  0;
		int_i[5] =  0;
		int_i[6] =  0;
		int_i[7] =  0;
		int_i[8] =  0;
		int_i[9] =  0;
		int_i[10] =  0;
		int_i[11] =  0;
		int_i[12] =  0;
		int_i[13] =  0;
		int_i[14] =  0;
		int_i[15] =  0;
		int_i[16] =  0;
		int_i[17] =  0;
		int_i[18] =  0;
		int_i[19] =  0;
		int_i[20] =  0;
		int_i[21] =  0;
		int_i[22] =  0;
		int_i[23] =  0;
		int_i[24] =  0;
		int_i[25] =  0;
		int_i[26] =  0;
		int_i[27] =  0;
		int_i[28] =  0;
		int_i[29] =  0;
		int_i[30] =  0;
		int_i[31] =  0;
		int_i[32] =  0;
		int_i[33] =  0;
		int_i[34] =  0;
		int_i[35] =  0;
		int_i[36] =  0;
		int_i[37] =  0;
		int_i[38] =  0;
		int_i[39] =  0;
		int_i[40] =  0;
		int_i[41] =  0;
		int_i[42] =  0;
		int_i[43] =  0;
		int_i[44] =  0;
		int_i[45] =  0;
		int_i[46] =  0;
		int_i[47] =  0;
		int_i[48] =  0;
		int_i[49] =  0;
		int_i[50] =  0;
		int_i[51] =  0;
		int_i[52] =  0;
		int_i[53] =  0;
		int_i[54] =  0;
		int_i[55] =  0;
		int_i[56] =  0;
		int_i[57] =  0;
		int_i[58] =  0;
		int_i[59] =  0;
		int_i[60] =  0;
		int_i[61] =  0;
		int_i[62] =  0;
		int_i[63] =  0;
		int_i[64] =  0;
		int_i[65] =  0;
		int_i[66] =  0;
		int_i[67] =  0;
		int_i[68] =  0;
		int_i[69] =  0;
		int_i[70] =  0;
		int_i[71] =  0;
		int_i[72] =  0;
		int_i[73] =  0;
		int_i[74] =  0;
		int_i[75] =  0;
		int_i[76] =  0;
		int_i[77] =  0;
		int_i[78] =  0;
		int_i[79] =  0;
		int_i[80] =  0;
		int_i[81] =  0;
		int_i[82] =  0;
		int_i[83] =  0;
		int_i[84] =  0;
		int_i[85] =  0;
		int_i[86] =  0;
		int_i[87] =  0;
		int_i[88] =  0;
		int_i[89] =  0;
		int_i[90] =  0;
		int_i[91] =  0;
		int_i[92] =  0;
		int_i[93] =  0;
		int_i[94] =  0;
		int_i[95] =  0;
		int_i[96] =  0;
		int_i[97] =  0;
		int_i[98] =  0;
		int_i[99] =  0;
		int_i[100] =  0;
		int_i[101] =  0;
		int_i[102] =  0;
		int_i[103] =  0;
		int_i[104] =  0;
		int_i[105] =  0;
		int_i[106] =  0;
		int_i[107] =  0;
		int_i[108] =  0;
		int_i[109] =  0;
		int_i[110] =  0;
		int_i[111] =  0;
		int_i[112] =  0;
		int_i[113] =  0;
		int_i[114] =  0;
		int_i[115] =  0;
		int_i[116] =  0;
		int_i[117] =  0;
		int_i[118] =  0;
		int_i[119] =  0;
		int_i[120] =  0;
		int_i[121] =  0;
		int_i[122] =  0;
		int_i[123] =  0;
		int_i[124] =  0;
		int_i[125] =  0;
		int_i[126] =  0;
		int_i[127] =  0;
		int_i[128] =  0;
		int_i[129] =  0;
		int_i[130] =  0;
		int_i[131] =  0;
		int_i[132] =  0;
		int_i[133] =  0;
		int_i[134] =  0;
		int_i[135] =  0;
		int_i[136] =  0;
		int_i[137] =  0;
		int_i[138] =  0;
		int_i[139] =  0;
		int_i[140] =  0;
		int_i[141] =  0;
		int_i[142] =  0;
		int_i[143] =  0;
		int_i[144] =  0;
		int_i[145] =  0;
		int_i[146] =  0;
		int_i[147] =  0;
		int_i[148] =  0;
		int_i[149] =  0;
		int_i[150] =  0;
		int_i[151] =  0;
		int_i[152] =  0;
		int_i[153] =  0;
		int_i[154] =  0;
		int_i[155] =  0;
		int_i[156] =  0;
		int_i[157] =  0;
		int_i[158] =  0;
		int_i[159] =  0;
		int_i[160] =  0;
		int_i[161] =  0;
		int_i[162] =  0;
		int_i[163] =  0;
		int_i[164] =  0;
		int_i[165] =  0;
		int_i[166] =  0;
		int_i[167] =  0;
		int_i[168] =  0;
		int_i[169] =  0;
		int_i[170] =  0;
		int_i[171] =  0;
		int_i[172] =  0;
		int_i[173] =  0;
		int_i[174] =  0;
		int_i[175] =  0;
		int_i[176] =  0;
		int_i[177] =  0;
		int_i[178] =  0;
		int_i[179] =  0;
		int_i[180] =  0;
		int_i[181] =  0;
		int_i[182] =  0;
		int_i[183] =  0;
		int_i[184] =  0;
		int_i[185] =  0;
		int_i[186] =  0;
		int_i[187] =  0;
		int_i[188] =  0;
		int_i[189] =  0;
		int_i[190] =  0;
		int_i[191] =  0;
		int_i[192] =  0;
		int_i[193] =  0;
		int_i[194] =  0;
		int_i[195] =  0;
		int_i[196] =  0;
		int_i[197] =  0;
		int_i[198] =  0;
		int_i[199] =  0;
		int_i[200] =  0;
		int_i[201] =  0;
		int_i[202] =  0;
		int_i[203] =  0;
		int_i[204] =  0;
		int_i[205] =  0;
		int_i[206] =  0;
		int_i[207] =  0;
		int_i[208] =  0;
		int_i[209] =  0;
		int_i[210] =  0;
		int_i[211] =  0;
		int_i[212] =  0;
		int_i[213] =  0;
		int_i[214] =  0;
		int_i[215] =  0;
		int_i[216] =  0;
		int_i[217] =  0;
		int_i[218] =  0;
		int_i[219] =  0;
		int_i[220] =  0;
		int_i[221] =  0;
		int_i[222] =  0;
		int_i[223] =  0;
		int_i[224] =  0;
		int_i[225] =  0;
		int_i[226] =  0;
		int_i[227] =  0;
		int_i[228] =  0;
		int_i[229] =  0;
		int_i[230] =  0;
		int_i[231] =  0;
		int_i[232] =  0;
		int_i[233] =  0;
		int_i[234] =  0;
		int_i[235] =  0;
		int_i[236] =  0;
		int_i[237] =  0;
		int_i[238] =  0;
		int_i[239] =  0;
		int_i[240] =  0;
		int_i[241] =  0;
		int_i[242] =  0;
		int_i[243] =  0;
		int_i[244] =  0;
		int_i[245] =  0;
		int_i[246] =  0;
		int_i[247] =  0;
		int_i[248] =  0;
		int_i[249] =  0;
		int_i[250] =  0;
		int_i[251] =  0;
		int_i[252] =  0;
		int_i[253] =  0;
		int_i[254] =  0;
		int_i[255] =  0;
		int_i[256] =  0;
		int_i[257] =  0;
		int_i[258] =  0;
		int_i[259] =  0;
		int_i[260] =  0;
		int_i[261] =  0;
		int_i[262] =  0;
		int_i[263] =  0;
		int_i[264] =  0;
		int_i[265] =  0;
		int_i[266] =  0;
		int_i[267] =  0;
		int_i[268] =  0;
		int_i[269] =  0;
		int_i[270] =  0;
		int_i[271] =  0;
		int_i[272] =  0;
		int_i[273] =  0;
		int_i[274] =  0;
		int_i[275] =  0;
		int_i[276] =  0;
		int_i[277] =  0;
		int_i[278] =  0;
		int_i[279] =  0;
		int_i[280] =  0;
		int_i[281] =  0;
		int_i[282] =  0;
		int_i[283] =  0;
		int_i[284] =  0;
		int_i[285] =  0;
		int_i[286] =  0;
		int_i[287] =  0;
		int_i[288] =  0;
		int_i[289] =  0;
		int_i[290] =  0;
		int_i[291] =  0;
		int_i[292] =  0;
		int_i[293] =  0;
		int_i[294] =  0;
		int_i[295] =  0;
		int_i[296] =  0;
		int_i[297] =  0;
		int_i[298] =  0;
		int_i[299] =  0;
		int_i[300] =  0;
		int_i[301] =  0;
		int_i[302] =  0;
		int_i[303] =  0;
		int_i[304] =  0;
		int_i[305] =  0;
		int_i[306] =  0;
		int_i[307] =  0;
		int_i[308] =  0;
		int_i[309] =  0;
		int_i[310] =  0;
		int_i[311] =  0;
		int_i[312] =  0;
		int_i[313] =  0;
		int_i[314] =  0;
		int_i[315] =  0;
		int_i[316] =  0;
		int_i[317] =  0;
		int_i[318] =  0;
		int_i[319] =  0;
		int_i[320] =  0;
		int_i[321] =  0;
		int_i[322] =  0;
		int_i[323] =  0;
		int_i[324] =  0;
		int_i[325] =  0;
		int_i[326] =  0;
		int_i[327] =  0;
		int_i[328] =  0;
		int_i[329] =  0;
		int_i[330] =  0;
		int_i[331] =  0;
		int_i[332] =  0;
		int_i[333] =  0;
		int_i[334] =  0;
		int_i[335] =  0;
		int_i[336] =  0;
		int_i[337] =  0;
		int_i[338] =  0;
		int_i[339] =  0;
		int_i[340] =  0;
		int_i[341] =  0;
		int_i[342] =  0;
		int_i[343] =  0;
		int_i[344] =  0;
		int_i[345] =  0;
		int_i[346] =  0;
		int_i[347] =  0;
		int_i[348] =  0;
		int_i[349] =  0;
		int_i[350] =  0;
		int_i[351] =  0;
		int_i[352] =  0;
		int_i[353] =  0;
		int_i[354] =  0;
		int_i[355] =  0;
		int_i[356] =  0;
		int_i[357] =  0;
		int_i[358] =  0;
		int_i[359] =  0;
		int_i[360] =  0;
		int_i[361] =  0;
		int_i[362] =  0;
		int_i[363] =  0;
		int_i[364] =  0;
		int_i[365] =  0;
		int_i[366] =  0;
		int_i[367] =  0;
		int_i[368] =  0;
		int_i[369] =  0;
		int_i[370] =  0;
		int_i[371] =  0;
		int_i[372] =  0;
		int_i[373] =  0;
		int_i[374] =  0;
		int_i[375] =  0;
		int_i[376] =  0;
		int_i[377] =  0;
		int_i[378] =  0;
		int_i[379] =  0;
		int_i[380] =  0;
		int_i[381] =  0;
		int_i[382] =  0;
		int_i[383] =  0;
		int_i[384] =  0;
		int_i[385] =  0;
		int_i[386] =  0;
		int_i[387] =  0;
		int_i[388] =  0;
		int_i[389] =  0;
		int_i[390] =  0;
		int_i[391] =  0;
		int_i[392] =  0;
		int_i[393] =  0;
		int_i[394] =  0;
		int_i[395] =  0;
		int_i[396] =  0;
		int_i[397] =  0;
		int_i[398] =  0;
		int_i[399] =  0;
		int_i[400] =  0;
		int_i[401] =  0;
		int_i[402] =  0;
		int_i[403] =  0;
		int_i[404] =  0;
		int_i[405] =  0;
		int_i[406] =  0;
		int_i[407] =  0;
		int_i[408] =  0;
		int_i[409] =  0;
		int_i[410] =  0;
		int_i[411] =  0;
		int_i[412] =  0;
		int_i[413] =  0;
		int_i[414] =  0;
		int_i[415] =  0;
		int_i[416] =  0;
		int_i[417] =  0;
		int_i[418] =  0;
		int_i[419] =  0;
		int_i[420] =  0;
		int_i[421] =  0;
		int_i[422] =  0;
		int_i[423] =  0;
		int_i[424] =  0;
		int_i[425] =  0;
		int_i[426] =  0;
		int_i[427] =  0;
		int_i[428] =  0;
		int_i[429] =  0;
		int_i[430] =  0;
		int_i[431] =  0;
		int_i[432] =  0;
		int_i[433] =  0;
		int_i[434] =  0;
		int_i[435] =  0;
		int_i[436] =  0;
		int_i[437] =  0;
		int_i[438] =  0;
		int_i[439] =  0;
		int_i[440] =  0;
		int_i[441] =  0;
		int_i[442] =  0;
		int_i[443] =  0;
		int_i[444] =  0;
		int_i[445] =  0;
		int_i[446] =  0;
		int_i[447] =  0;
		int_i[448] =  0;
		int_i[449] =  0;
		int_i[450] =  0;
		int_i[451] =  0;
		int_i[452] =  0;
		int_i[453] =  0;
		int_i[454] =  0;
		int_i[455] =  0;
		int_i[456] =  0;
		int_i[457] =  0;
		int_i[458] =  0;
		int_i[459] =  0;
		int_i[460] =  0;
		int_i[461] =  0;
		int_i[462] =  0;
		int_i[463] =  0;
		int_i[464] =  0;
		int_i[465] =  0;
		int_i[466] =  0;
		int_i[467] =  0;
		int_i[468] =  0;
		int_i[469] =  0;
		int_i[470] =  0;
		int_i[471] =  0;
		int_i[472] =  0;
		int_i[473] =  0;
		int_i[474] =  0;
		int_i[475] =  0;
		int_i[476] =  0;
		int_i[477] =  0;
		int_i[478] =  0;
		int_i[479] =  0;
		int_i[480] =  0;
		int_i[481] =  0;
		int_i[482] =  0;
		int_i[483] =  0;
		int_i[484] =  0;
		int_i[485] =  0;
		int_i[486] =  0;
		int_i[487] =  0;
		int_i[488] =  0;
		int_i[489] =  0;
		int_i[490] =  0;
		int_i[491] =  0;
		int_i[492] =  0;
		int_i[493] =  0;
		int_i[494] =  0;
		int_i[495] =  0;
		int_i[496] =  0;
		int_i[497] =  0;
		int_i[498] =  0;
		int_i[499] =  0;
		int_i[500] =  0;
		int_i[501] =  0;
		int_i[502] =  0;
		int_i[503] =  0;
		int_i[504] =  0;
		int_i[505] =  0;
		int_i[506] =  0;
		int_i[507] =  0;
		int_i[508] =  0;
		int_i[509] =  0;
		int_i[510] =  0;
		int_i[511] =  0;
		int_i[512] =  0;
		int_i[513] =  0;
		int_i[514] =  0;
		int_i[515] =  0;
		int_i[516] =  0;
		int_i[517] =  0;
		int_i[518] =  0;
		int_i[519] =  0;
		int_i[520] =  0;
		int_i[521] =  0;
		int_i[522] =  0;
		int_i[523] =  0;
		int_i[524] =  0;
		int_i[525] =  0;
		int_i[526] =  0;
		int_i[527] =  0;
		int_i[528] =  0;
		int_i[529] =  0;
		int_i[530] =  0;
		int_i[531] =  0;
		int_i[532] =  0;
		int_i[533] =  0;
		int_i[534] =  0;
		int_i[535] =  0;
		int_i[536] =  0;
		int_i[537] =  0;
		int_i[538] =  0;
		int_i[539] =  0;
		int_i[540] =  0;
		int_i[541] =  0;
		int_i[542] =  0;
		int_i[543] =  0;
		int_i[544] =  0;
		int_i[545] =  0;
		int_i[546] =  0;
		int_i[547] =  0;
		int_i[548] =  0;
		int_i[549] =  0;
		int_i[550] =  0;
		int_i[551] =  0;
		int_i[552] =  0;
		int_i[553] =  0;
		int_i[554] =  0;
		int_i[555] =  0;
		int_i[556] =  0;
		int_i[557] =  0;
		int_i[558] =  0;
		int_i[559] =  0;
		int_i[560] =  0;
		int_i[561] =  0;
		int_i[562] =  0;
		int_i[563] =  0;
		int_i[564] =  0;
		int_i[565] =  0;
		int_i[566] =  0;
		int_i[567] =  0;
		int_i[568] =  0;
		int_i[569] =  0;
		int_i[570] =  0;
		int_i[571] =  0;
		int_i[572] =  0;
		int_i[573] =  0;
		int_i[574] =  0;
		int_i[575] =  0;
		int_i[576] =  0;
		int_i[577] =  0;
		int_i[578] =  0;
		int_i[579] =  0;
		int_i[580] =  0;
		int_i[581] =  0;
		int_i[582] =  0;
		int_i[583] =  0;
		int_i[584] =  0;
		int_i[585] =  0;
		int_i[586] =  0;
		int_i[587] =  0;
		int_i[588] =  0;
		int_i[589] =  0;
		int_i[590] =  0;
		int_i[591] =  0;
		int_i[592] =  0;
		int_i[593] =  0;
		int_i[594] =  0;
		int_i[595] =  0;
		int_i[596] =  0;
		int_i[597] =  0;
		int_i[598] =  0;
		int_i[599] =  0;
		int_i[600] =  0;
		int_i[601] =  0;
		int_i[602] =  0;
		int_i[603] =  0;
		int_i[604] =  0;
		int_i[605] =  0;
		int_i[606] =  0;
		int_i[607] =  0;
		int_i[608] =  0;
		int_i[609] =  0;
		int_i[610] =  0;
		int_i[611] =  0;
		int_i[612] =  0;
		int_i[613] =  0;
		int_i[614] =  0;
		int_i[615] =  0;
		int_i[616] =  0;
		int_i[617] =  0;
		int_i[618] =  0;
		int_i[619] =  0;
		int_i[620] =  0;
		int_i[621] =  0;
		int_i[622] =  0;
		int_i[623] =  0;
		int_i[624] =  0;
		int_i[625] =  0;
		int_i[626] =  0;
		int_i[627] =  0;
		int_i[628] =  0;
		int_i[629] =  0;
		int_i[630] =  0;
		int_i[631] =  0;
		int_i[632] =  0;
		int_i[633] =  0;
		int_i[634] =  0;
		int_i[635] =  0;
		int_i[636] =  0;
		int_i[637] =  0;
		int_i[638] =  0;
		int_i[639] =  0;
		int_i[640] =  0;
		int_i[641] =  0;
		int_i[642] =  0;
		int_i[643] =  0;
		int_i[644] =  0;
		int_i[645] =  0;
		int_i[646] =  0;
		int_i[647] =  0;
		int_i[648] =  0;
		int_i[649] =  0;
		int_i[650] =  0;
		int_i[651] =  0;
		int_i[652] =  0;
		int_i[653] =  0;
		int_i[654] =  0;
		int_i[655] =  0;
		int_i[656] =  0;
		int_i[657] =  0;
		int_i[658] =  0;
		int_i[659] =  0;
		int_i[660] =  0;
		int_i[661] =  0;
		int_i[662] =  0;
		int_i[663] =  0;
		int_i[664] =  0;
		int_i[665] =  0;
		int_i[666] =  0;
		int_i[667] =  0;
		int_i[668] =  0;
		int_i[669] =  0;
		int_i[670] =  0;
		int_i[671] =  0;
		int_i[672] =  0;
		int_i[673] =  0;
		int_i[674] =  0;
		int_i[675] =  0;
		int_i[676] =  0;
		int_i[677] =  0;
		int_i[678] =  0;
		int_i[679] =  0;
		int_i[680] =  0;
		int_i[681] =  0;
		int_i[682] =  0;
		int_i[683] =  0;
		int_i[684] =  0;
		int_i[685] =  0;
		int_i[686] =  0;
		int_i[687] =  0;
		int_i[688] =  0;
		int_i[689] =  0;
		int_i[690] =  0;
		int_i[691] =  0;
		int_i[692] =  0;
		int_i[693] =  0;
		int_i[694] =  0;
		int_i[695] =  0;
		int_i[696] =  0;
		int_i[697] =  0;
		int_i[698] =  0;
		int_i[699] =  0;
		int_i[700] =  0;
		int_i[701] =  0;
		int_i[702] =  0;
		int_i[703] =  0;
		int_i[704] =  0;
		int_i[705] =  0;
		int_i[706] =  0;
		int_i[707] =  0;
		int_i[708] =  0;
		int_i[709] =  0;
		int_i[710] =  0;
		int_i[711] =  0;
		int_i[712] =  0;
		int_i[713] =  0;
		int_i[714] =  0;
		int_i[715] =  0;
		int_i[716] =  0;
		int_i[717] =  0;
		int_i[718] =  0;
		int_i[719] =  0;
		int_i[720] =  0;
		int_i[721] =  0;
		int_i[722] =  0;
		int_i[723] =  0;
		int_i[724] =  0;
		int_i[725] =  0;
		int_i[726] =  0;
		int_i[727] =  0;
		int_i[728] =  0;
		int_i[729] =  0;
		int_i[730] =  0;
		int_i[731] =  0;
		int_i[732] =  0;
		int_i[733] =  0;
		int_i[734] =  0;
		int_i[735] =  0;
		int_i[736] =  0;
		int_i[737] =  0;
		int_i[738] =  0;
		int_i[739] =  0;
		int_i[740] =  0;
		int_i[741] =  0;
		int_i[742] =  0;
		int_i[743] =  0;
		int_i[744] =  0;
		int_i[745] =  0;
		int_i[746] =  0;
		int_i[747] =  0;
		int_i[748] =  0;
		int_i[749] =  0;
		int_i[750] =  0;
		int_i[751] =  0;
		int_i[752] =  0;
		int_i[753] =  0;
		int_i[754] =  0;
		int_i[755] =  0;
		int_i[756] =  0;
		int_i[757] =  0;
		int_i[758] =  0;
		int_i[759] =  0;
		int_i[760] =  0;
		int_i[761] =  0;
		int_i[762] =  0;
		int_i[763] =  0;
		int_i[764] =  0;
		int_i[765] =  0;
		int_i[766] =  0;
		int_i[767] =  0;
		int_i[768] =  0;
		int_i[769] =  0;
		int_i[770] =  0;
		int_i[771] =  0;
		int_i[772] =  0;
		int_i[773] =  0;
		int_i[774] =  0;
		int_i[775] =  0;
		int_i[776] =  0;
		int_i[777] =  0;
		int_i[778] =  0;
		int_i[779] =  0;
		int_i[780] =  0;
		int_i[781] =  0;
		int_i[782] =  0;
		int_i[783] =  0;
		int_i[784] =  0;
		int_i[785] =  0;
		int_i[786] =  0;
		int_i[787] =  0;
		int_i[788] =  0;
		int_i[789] =  0;
		int_i[790] =  0;
		int_i[791] =  0;
		int_i[792] =  0;
		int_i[793] =  0;
		int_i[794] =  0;
		int_i[795] =  0;
		int_i[796] =  0;
		int_i[797] =  0;
		int_i[798] =  0;
		int_i[799] =  0;
		int_i[800] =  0;
		int_i[801] =  0;
		int_i[802] =  0;
		int_i[803] =  0;
		int_i[804] =  0;
		int_i[805] =  0;
		int_i[806] =  0;
		int_i[807] =  0;
		int_i[808] =  0;
		int_i[809] =  0;
		int_i[810] =  0;
		int_i[811] =  0;
		int_i[812] =  0;
		int_i[813] =  0;
		int_i[814] =  0;
		int_i[815] =  0;
		int_i[816] =  0;
		int_i[817] =  0;
		int_i[818] =  0;
		int_i[819] =  0;
		int_i[820] =  0;
		int_i[821] =  0;
		int_i[822] =  0;
		int_i[823] =  0;
		int_i[824] =  0;
		int_i[825] =  0;
		int_i[826] =  0;
		int_i[827] =  0;
		int_i[828] =  0;
		int_i[829] =  0;
		int_i[830] =  0;
		int_i[831] =  0;
		int_i[832] =  0;
		int_i[833] =  0;
		int_i[834] =  0;
		int_i[835] =  0;
		int_i[836] =  0;
		int_i[837] =  0;
		int_i[838] =  0;
		int_i[839] =  0;
		int_i[840] =  0;
		int_i[841] =  0;
		int_i[842] =  0;
		int_i[843] =  0;
		int_i[844] =  0;
		int_i[845] =  0;
		int_i[846] =  0;
		int_i[847] =  0;
		int_i[848] =  0;
		int_i[849] =  0;
		int_i[850] =  0;
		int_i[851] =  0;
		int_i[852] =  0;
		int_i[853] =  0;
		int_i[854] =  0;
		int_i[855] =  0;
		int_i[856] =  0;
		int_i[857] =  0;
		int_i[858] =  0;
		int_i[859] =  0;
		int_i[860] =  0;
		int_i[861] =  0;
		int_i[862] =  0;
		int_i[863] =  0;
		int_i[864] =  0;
		int_i[865] =  0;
		int_i[866] =  0;
		int_i[867] =  0;
		int_i[868] =  0;
		int_i[869] =  0;
		int_i[870] =  0;
		int_i[871] =  0;
		int_i[872] =  0;
		int_i[873] =  0;
		int_i[874] =  0;
		int_i[875] =  0;
		int_i[876] =  0;
		int_i[877] =  0;
		int_i[878] =  0;
		int_i[879] =  0;
		int_i[880] =  0;
		int_i[881] =  0;
		int_i[882] =  0;
		int_i[883] =  0;
		int_i[884] =  0;
		int_i[885] =  0;
		int_i[886] =  0;
		int_i[887] =  0;
		int_i[888] =  0;
		int_i[889] =  0;
		int_i[890] =  0;
		int_i[891] =  0;
		int_i[892] =  0;
		int_i[893] =  0;
		int_i[894] =  0;
		int_i[895] =  0;
		int_i[896] =  0;
		int_i[897] =  0;
		int_i[898] =  0;
		int_i[899] =  0;
		int_i[900] =  0;
		int_i[901] =  0;
		int_i[902] =  0;
		int_i[903] =  0;
		int_i[904] =  0;
		int_i[905] =  0;
		int_i[906] =  0;
		int_i[907] =  0;
		int_i[908] =  0;
		int_i[909] =  0;
		int_i[910] =  0;
		int_i[911] =  0;
		int_i[912] =  0;
		int_i[913] =  0;
		int_i[914] =  0;
		int_i[915] =  0;
		int_i[916] =  0;
		int_i[917] =  0;
		int_i[918] =  0;
		int_i[919] =  0;
		int_i[920] =  0;
		int_i[921] =  0;
		int_i[922] =  0;
		int_i[923] =  0;
		int_i[924] =  0;
		int_i[925] =  0;
		int_i[926] =  0;
		int_i[927] =  0;
		int_i[928] =  0;
		int_i[929] =  0;
		int_i[930] =  0;
		int_i[931] =  0;
		int_i[932] =  0;
		int_i[933] =  0;
		int_i[934] =  0;
		int_i[935] =  0;
		int_i[936] =  0;
		int_i[937] =  0;
		int_i[938] =  0;
		int_i[939] =  0;
		int_i[940] =  0;
		int_i[941] =  0;
		int_i[942] =  0;
		int_i[943] =  0;
		int_i[944] =  0;
		int_i[945] =  0;
		int_i[946] =  0;
		int_i[947] =  0;
		int_i[948] =  0;
		int_i[949] =  0;
		int_i[950] =  0;
		int_i[951] =  0;
		int_i[952] =  0;
		int_i[953] =  0;
		int_i[954] =  0;
		int_i[955] =  0;
		int_i[956] =  0;
		int_i[957] =  0;
		int_i[958] =  0;
		int_i[959] =  0;
		int_i[960] =  0;
		int_i[961] =  0;
		int_i[962] =  0;
		int_i[963] =  0;
		int_i[964] =  0;
		int_i[965] =  0;
		int_i[966] =  0;
		int_i[967] =  0;
		int_i[968] =  0;
		int_i[969] =  0;
		int_i[970] =  0;
		int_i[971] =  0;
		int_i[972] =  0;
		int_i[973] =  0;
		int_i[974] =  0;
		int_i[975] =  0;
		int_i[976] =  0;
		int_i[977] =  0;
		int_i[978] =  0;
		int_i[979] =  0;
		int_i[980] =  0;
		int_i[981] =  0;
		int_i[982] =  0;
		int_i[983] =  0;
		int_i[984] =  0;
		int_i[985] =  0;
		int_i[986] =  0;
		int_i[987] =  0;
		int_i[988] =  0;
		int_i[989] =  0;
		int_i[990] =  0;
		int_i[991] =  0;
		int_i[992] =  0;
		int_i[993] =  0;
		int_i[994] =  0;
		int_i[995] =  0;
		int_i[996] =  0;
		int_i[997] =  0;
		int_i[998] =  0;
		int_i[999] =  0;
		int_i[1000] =  0;
		int_i[1001] =  0;
		int_i[1002] =  0;
		int_i[1003] =  0;
		int_i[1004] =  0;
		int_i[1005] =  0;
		int_i[1006] =  0;
		int_i[1007] =  0;
		int_i[1008] =  0;
		int_i[1009] =  0;
		int_i[1010] =  0;
		int_i[1011] =  0;
		int_i[1012] =  0;
		int_i[1013] =  0;
		int_i[1014] =  0;
		int_i[1015] =  0;
		int_i[1016] =  0;
		int_i[1017] =  0;
		int_i[1018] =  0;
		int_i[1019] =  0;
		int_i[1020] =  0;
		int_i[1021] =  0;
		int_i[1022] =  0;
		int_i[1023] =  0;
	end
////////////////////////////////////////////	
	initial begin
		clk       = 0;
		rst_n     = 1;
		in_valid  = 0;
		@(negedge clk);
		@(negedge clk) rst_n = 0;
		@(negedge clk) rst_n = 1;
		@(negedge clk);
		////////////////////////
		for(j=0;j<FFT_size;j=j+1) begin
			@(negedge clk);
			in_valid 	= 1;
			din_r 		= int_r[j];
			din_i 		= int_i[j];
		end
		@(negedge clk) in_valid = 0;		
		////////////////////////
		////////////////////////		
		for(j=0;j<FFT_size;j=j+1) begin
			while(!out_valid) begin
				@(negedge clk); 
			end	
			@(negedge clk);
		end
		///////////////////////
		///////////////////////		
		$stop;
	end
endmodule
